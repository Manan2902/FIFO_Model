// This is the unpowered netlist.
module FIFO_Model (Clk,
    FClrN,
    FInN,
    FOutN,
    F_EmptyN,
    F_FirstN,
    F_FullN,
    F_LastN,
    F_SLastN,
    RstN,
    Data_In,
    F_Data);
 input Clk;
 input FClrN;
 input FInN;
 input FOutN;
 output F_EmptyN;
 output F_FirstN;
 output F_FullN;
 output F_LastN;
 output F_SLastN;
 input RstN;
 input [31:0] Data_In;
 output [31:0] F_Data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire clknet_0_Clk;
 wire clknet_4_0_0_Clk;
 wire clknet_4_10_0_Clk;
 wire clknet_4_11_0_Clk;
 wire clknet_4_12_0_Clk;
 wire clknet_4_13_0_Clk;
 wire clknet_4_14_0_Clk;
 wire clknet_4_15_0_Clk;
 wire clknet_4_1_0_Clk;
 wire clknet_4_2_0_Clk;
 wire clknet_4_3_0_Clk;
 wire clknet_4_4_0_Clk;
 wire clknet_4_5_0_Clk;
 wire clknet_4_6_0_Clk;
 wire clknet_4_7_0_Clk;
 wire clknet_4_8_0_Clk;
 wire clknet_4_9_0_Clk;
 wire \fcounter[0] ;
 wire \fcounter[1] ;
 wire \fcounter[2] ;
 wire \memblk.FIFO[0][0] ;
 wire \memblk.FIFO[0][10] ;
 wire \memblk.FIFO[0][11] ;
 wire \memblk.FIFO[0][12] ;
 wire \memblk.FIFO[0][13] ;
 wire \memblk.FIFO[0][14] ;
 wire \memblk.FIFO[0][15] ;
 wire \memblk.FIFO[0][16] ;
 wire \memblk.FIFO[0][17] ;
 wire \memblk.FIFO[0][18] ;
 wire \memblk.FIFO[0][19] ;
 wire \memblk.FIFO[0][1] ;
 wire \memblk.FIFO[0][20] ;
 wire \memblk.FIFO[0][21] ;
 wire \memblk.FIFO[0][22] ;
 wire \memblk.FIFO[0][23] ;
 wire \memblk.FIFO[0][24] ;
 wire \memblk.FIFO[0][25] ;
 wire \memblk.FIFO[0][26] ;
 wire \memblk.FIFO[0][27] ;
 wire \memblk.FIFO[0][28] ;
 wire \memblk.FIFO[0][29] ;
 wire \memblk.FIFO[0][2] ;
 wire \memblk.FIFO[0][30] ;
 wire \memblk.FIFO[0][31] ;
 wire \memblk.FIFO[0][3] ;
 wire \memblk.FIFO[0][4] ;
 wire \memblk.FIFO[0][5] ;
 wire \memblk.FIFO[0][6] ;
 wire \memblk.FIFO[0][7] ;
 wire \memblk.FIFO[0][8] ;
 wire \memblk.FIFO[0][9] ;
 wire \memblk.FIFO[1][0] ;
 wire \memblk.FIFO[1][10] ;
 wire \memblk.FIFO[1][11] ;
 wire \memblk.FIFO[1][12] ;
 wire \memblk.FIFO[1][13] ;
 wire \memblk.FIFO[1][14] ;
 wire \memblk.FIFO[1][15] ;
 wire \memblk.FIFO[1][16] ;
 wire \memblk.FIFO[1][17] ;
 wire \memblk.FIFO[1][18] ;
 wire \memblk.FIFO[1][19] ;
 wire \memblk.FIFO[1][1] ;
 wire \memblk.FIFO[1][20] ;
 wire \memblk.FIFO[1][21] ;
 wire \memblk.FIFO[1][22] ;
 wire \memblk.FIFO[1][23] ;
 wire \memblk.FIFO[1][24] ;
 wire \memblk.FIFO[1][25] ;
 wire \memblk.FIFO[1][26] ;
 wire \memblk.FIFO[1][27] ;
 wire \memblk.FIFO[1][28] ;
 wire \memblk.FIFO[1][29] ;
 wire \memblk.FIFO[1][2] ;
 wire \memblk.FIFO[1][30] ;
 wire \memblk.FIFO[1][31] ;
 wire \memblk.FIFO[1][3] ;
 wire \memblk.FIFO[1][4] ;
 wire \memblk.FIFO[1][5] ;
 wire \memblk.FIFO[1][6] ;
 wire \memblk.FIFO[1][7] ;
 wire \memblk.FIFO[1][8] ;
 wire \memblk.FIFO[1][9] ;
 wire \memblk.FIFO[2][0] ;
 wire \memblk.FIFO[2][10] ;
 wire \memblk.FIFO[2][11] ;
 wire \memblk.FIFO[2][12] ;
 wire \memblk.FIFO[2][13] ;
 wire \memblk.FIFO[2][14] ;
 wire \memblk.FIFO[2][15] ;
 wire \memblk.FIFO[2][16] ;
 wire \memblk.FIFO[2][17] ;
 wire \memblk.FIFO[2][18] ;
 wire \memblk.FIFO[2][19] ;
 wire \memblk.FIFO[2][1] ;
 wire \memblk.FIFO[2][20] ;
 wire \memblk.FIFO[2][21] ;
 wire \memblk.FIFO[2][22] ;
 wire \memblk.FIFO[2][23] ;
 wire \memblk.FIFO[2][24] ;
 wire \memblk.FIFO[2][25] ;
 wire \memblk.FIFO[2][26] ;
 wire \memblk.FIFO[2][27] ;
 wire \memblk.FIFO[2][28] ;
 wire \memblk.FIFO[2][29] ;
 wire \memblk.FIFO[2][2] ;
 wire \memblk.FIFO[2][30] ;
 wire \memblk.FIFO[2][31] ;
 wire \memblk.FIFO[2][3] ;
 wire \memblk.FIFO[2][4] ;
 wire \memblk.FIFO[2][5] ;
 wire \memblk.FIFO[2][6] ;
 wire \memblk.FIFO[2][7] ;
 wire \memblk.FIFO[2][8] ;
 wire \memblk.FIFO[2][9] ;
 wire \memblk.FIFO[3][0] ;
 wire \memblk.FIFO[3][10] ;
 wire \memblk.FIFO[3][11] ;
 wire \memblk.FIFO[3][12] ;
 wire \memblk.FIFO[3][13] ;
 wire \memblk.FIFO[3][14] ;
 wire \memblk.FIFO[3][15] ;
 wire \memblk.FIFO[3][16] ;
 wire \memblk.FIFO[3][17] ;
 wire \memblk.FIFO[3][18] ;
 wire \memblk.FIFO[3][19] ;
 wire \memblk.FIFO[3][1] ;
 wire \memblk.FIFO[3][20] ;
 wire \memblk.FIFO[3][21] ;
 wire \memblk.FIFO[3][22] ;
 wire \memblk.FIFO[3][23] ;
 wire \memblk.FIFO[3][24] ;
 wire \memblk.FIFO[3][25] ;
 wire \memblk.FIFO[3][26] ;
 wire \memblk.FIFO[3][27] ;
 wire \memblk.FIFO[3][28] ;
 wire \memblk.FIFO[3][29] ;
 wire \memblk.FIFO[3][2] ;
 wire \memblk.FIFO[3][30] ;
 wire \memblk.FIFO[3][31] ;
 wire \memblk.FIFO[3][3] ;
 wire \memblk.FIFO[3][4] ;
 wire \memblk.FIFO[3][5] ;
 wire \memblk.FIFO[3][6] ;
 wire \memblk.FIFO[3][7] ;
 wire \memblk.FIFO[3][8] ;
 wire \memblk.FIFO[3][9] ;
 wire \memblk.rd_addr[0] ;
 wire \memblk.rd_addr[1] ;
 wire \memblk.wr_addr[0] ;
 wire \memblk.wr_addr[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_127 ();
 sky130_fd_sc_hd__clkbuf_2 _389_ (.A(\memblk.rd_addr[0] ),
    .X(_140_));
 sky130_fd_sc_hd__buf_2 _390_ (.A(_140_),
    .X(_141_));
 sky130_fd_sc_hd__clkbuf_2 _391_ (.A(\memblk.rd_addr[1] ),
    .X(_142_));
 sky130_fd_sc_hd__clkbuf_2 _392_ (.A(_142_),
    .X(_143_));
 sky130_fd_sc_hd__mux4_1 _393_ (.A0(\memblk.FIFO[0][0] ),
    .A1(\memblk.FIFO[1][0] ),
    .A2(\memblk.FIFO[2][0] ),
    .A3(\memblk.FIFO[3][0] ),
    .S0(_141_),
    .S1(_143_),
    .X(_144_));
 sky130_fd_sc_hd__clkbuf_1 _394_ (.A(_144_),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 _395_ (.A0(\memblk.FIFO[0][1] ),
    .A1(\memblk.FIFO[1][1] ),
    .A2(\memblk.FIFO[2][1] ),
    .A3(\memblk.FIFO[3][1] ),
    .S0(_141_),
    .S1(_143_),
    .X(_145_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(_145_),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 _397_ (.A0(\memblk.FIFO[0][2] ),
    .A1(\memblk.FIFO[1][2] ),
    .A2(\memblk.FIFO[2][2] ),
    .A3(\memblk.FIFO[3][2] ),
    .S0(_141_),
    .S1(_143_),
    .X(_146_));
 sky130_fd_sc_hd__clkbuf_1 _398_ (.A(_146_),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 _399_ (.A0(\memblk.FIFO[0][3] ),
    .A1(\memblk.FIFO[1][3] ),
    .A2(\memblk.FIFO[2][3] ),
    .A3(\memblk.FIFO[3][3] ),
    .S0(_141_),
    .S1(_143_),
    .X(_147_));
 sky130_fd_sc_hd__clkbuf_1 _400_ (.A(_147_),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 _401_ (.A0(\memblk.FIFO[0][4] ),
    .A1(\memblk.FIFO[1][4] ),
    .A2(\memblk.FIFO[2][4] ),
    .A3(\memblk.FIFO[3][4] ),
    .S0(_141_),
    .S1(_143_),
    .X(_148_));
 sky130_fd_sc_hd__clkbuf_1 _402_ (.A(_148_),
    .X(net63));
 sky130_fd_sc_hd__buf_2 _403_ (.A(_140_),
    .X(_149_));
 sky130_fd_sc_hd__clkbuf_2 _404_ (.A(_142_),
    .X(_150_));
 sky130_fd_sc_hd__mux4_1 _405_ (.A0(\memblk.FIFO[0][5] ),
    .A1(\memblk.FIFO[1][5] ),
    .A2(\memblk.FIFO[2][5] ),
    .A3(\memblk.FIFO[3][5] ),
    .S0(_149_),
    .S1(_150_),
    .X(_151_));
 sky130_fd_sc_hd__clkbuf_1 _406_ (.A(_151_),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 _407_ (.A0(\memblk.FIFO[0][6] ),
    .A1(\memblk.FIFO[1][6] ),
    .A2(\memblk.FIFO[2][6] ),
    .A3(\memblk.FIFO[3][6] ),
    .S0(_149_),
    .S1(_150_),
    .X(_152_));
 sky130_fd_sc_hd__clkbuf_1 _408_ (.A(_152_),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 _409_ (.A0(\memblk.FIFO[0][7] ),
    .A1(\memblk.FIFO[1][7] ),
    .A2(\memblk.FIFO[2][7] ),
    .A3(\memblk.FIFO[3][7] ),
    .S0(_149_),
    .S1(_150_),
    .X(_153_));
 sky130_fd_sc_hd__clkbuf_1 _410_ (.A(_153_),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 _411_ (.A0(\memblk.FIFO[0][8] ),
    .A1(\memblk.FIFO[1][8] ),
    .A2(\memblk.FIFO[2][8] ),
    .A3(\memblk.FIFO[3][8] ),
    .S0(_149_),
    .S1(_150_),
    .X(_154_));
 sky130_fd_sc_hd__clkbuf_1 _412_ (.A(_154_),
    .X(net67));
 sky130_fd_sc_hd__mux4_1 _413_ (.A0(\memblk.FIFO[0][9] ),
    .A1(\memblk.FIFO[1][9] ),
    .A2(\memblk.FIFO[2][9] ),
    .A3(\memblk.FIFO[3][9] ),
    .S0(_149_),
    .S1(_150_),
    .X(_155_));
 sky130_fd_sc_hd__clkbuf_1 _414_ (.A(_155_),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 _415_ (.A0(\memblk.FIFO[0][10] ),
    .A1(\memblk.FIFO[1][10] ),
    .A2(\memblk.FIFO[2][10] ),
    .A3(\memblk.FIFO[3][10] ),
    .S0(_149_),
    .S1(_150_),
    .X(_156_));
 sky130_fd_sc_hd__clkbuf_1 _416_ (.A(_156_),
    .X(net38));
 sky130_fd_sc_hd__buf_2 _417_ (.A(\memblk.rd_addr[0] ),
    .X(_157_));
 sky130_fd_sc_hd__clkbuf_2 _418_ (.A(_142_),
    .X(_158_));
 sky130_fd_sc_hd__mux4_1 _419_ (.A0(\memblk.FIFO[0][11] ),
    .A1(\memblk.FIFO[1][11] ),
    .A2(\memblk.FIFO[2][11] ),
    .A3(\memblk.FIFO[3][11] ),
    .S0(_157_),
    .S1(_158_),
    .X(_159_));
 sky130_fd_sc_hd__clkbuf_1 _420_ (.A(_159_),
    .X(net39));
 sky130_fd_sc_hd__mux4_1 _421_ (.A0(\memblk.FIFO[0][12] ),
    .A1(\memblk.FIFO[1][12] ),
    .A2(\memblk.FIFO[2][12] ),
    .A3(\memblk.FIFO[3][12] ),
    .S0(_157_),
    .S1(_158_),
    .X(_160_));
 sky130_fd_sc_hd__clkbuf_1 _422_ (.A(_160_),
    .X(net40));
 sky130_fd_sc_hd__mux4_1 _423_ (.A0(\memblk.FIFO[0][13] ),
    .A1(\memblk.FIFO[1][13] ),
    .A2(\memblk.FIFO[2][13] ),
    .A3(\memblk.FIFO[3][13] ),
    .S0(_157_),
    .S1(_158_),
    .X(_161_));
 sky130_fd_sc_hd__clkbuf_1 _424_ (.A(_161_),
    .X(net41));
 sky130_fd_sc_hd__mux4_1 _425_ (.A0(\memblk.FIFO[0][14] ),
    .A1(\memblk.FIFO[1][14] ),
    .A2(\memblk.FIFO[2][14] ),
    .A3(\memblk.FIFO[3][14] ),
    .S0(_157_),
    .S1(_158_),
    .X(_162_));
 sky130_fd_sc_hd__clkbuf_1 _426_ (.A(_162_),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 _427_ (.A0(\memblk.FIFO[0][15] ),
    .A1(\memblk.FIFO[1][15] ),
    .A2(\memblk.FIFO[2][15] ),
    .A3(\memblk.FIFO[3][15] ),
    .S0(_157_),
    .S1(_158_),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_1 _428_ (.A(_163_),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 _429_ (.A0(\memblk.FIFO[0][16] ),
    .A1(\memblk.FIFO[1][16] ),
    .A2(\memblk.FIFO[2][16] ),
    .A3(\memblk.FIFO[3][16] ),
    .S0(_157_),
    .S1(_158_),
    .X(_164_));
 sky130_fd_sc_hd__clkbuf_1 _430_ (.A(_164_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 _431_ (.A(\memblk.rd_addr[0] ),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_2 _432_ (.A(\memblk.rd_addr[1] ),
    .X(_166_));
 sky130_fd_sc_hd__mux4_1 _433_ (.A0(\memblk.FIFO[0][17] ),
    .A1(\memblk.FIFO[1][17] ),
    .A2(\memblk.FIFO[2][17] ),
    .A3(\memblk.FIFO[3][17] ),
    .S0(_165_),
    .S1(_166_),
    .X(_167_));
 sky130_fd_sc_hd__clkbuf_1 _434_ (.A(_167_),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 _435_ (.A0(\memblk.FIFO[0][18] ),
    .A1(\memblk.FIFO[1][18] ),
    .A2(\memblk.FIFO[2][18] ),
    .A3(\memblk.FIFO[3][18] ),
    .S0(_165_),
    .S1(_166_),
    .X(_168_));
 sky130_fd_sc_hd__clkbuf_1 _436_ (.A(_168_),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 _437_ (.A0(\memblk.FIFO[0][19] ),
    .A1(\memblk.FIFO[1][19] ),
    .A2(\memblk.FIFO[2][19] ),
    .A3(\memblk.FIFO[3][19] ),
    .S0(_165_),
    .S1(_166_),
    .X(_169_));
 sky130_fd_sc_hd__clkbuf_1 _438_ (.A(_169_),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 _439_ (.A0(\memblk.FIFO[0][20] ),
    .A1(\memblk.FIFO[1][20] ),
    .A2(\memblk.FIFO[2][20] ),
    .A3(\memblk.FIFO[3][20] ),
    .S0(_165_),
    .S1(_166_),
    .X(_170_));
 sky130_fd_sc_hd__clkbuf_1 _440_ (.A(_170_),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 _441_ (.A0(\memblk.FIFO[0][21] ),
    .A1(\memblk.FIFO[1][21] ),
    .A2(\memblk.FIFO[2][21] ),
    .A3(\memblk.FIFO[3][21] ),
    .S0(_165_),
    .S1(_166_),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _442_ (.A(_171_),
    .X(net50));
 sky130_fd_sc_hd__mux4_1 _443_ (.A0(\memblk.FIFO[0][22] ),
    .A1(\memblk.FIFO[1][22] ),
    .A2(\memblk.FIFO[2][22] ),
    .A3(\memblk.FIFO[3][22] ),
    .S0(_165_),
    .S1(_166_),
    .X(_172_));
 sky130_fd_sc_hd__clkbuf_1 _444_ (.A(_172_),
    .X(net51));
 sky130_fd_sc_hd__buf_2 _445_ (.A(\memblk.rd_addr[0] ),
    .X(_173_));
 sky130_fd_sc_hd__clkbuf_2 _446_ (.A(\memblk.rd_addr[1] ),
    .X(_174_));
 sky130_fd_sc_hd__mux4_1 _447_ (.A0(\memblk.FIFO[0][23] ),
    .A1(\memblk.FIFO[1][23] ),
    .A2(\memblk.FIFO[2][23] ),
    .A3(\memblk.FIFO[3][23] ),
    .S0(_173_),
    .S1(_174_),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_1 _448_ (.A(_175_),
    .X(net52));
 sky130_fd_sc_hd__mux4_1 _449_ (.A0(\memblk.FIFO[0][24] ),
    .A1(\memblk.FIFO[1][24] ),
    .A2(\memblk.FIFO[2][24] ),
    .A3(\memblk.FIFO[3][24] ),
    .S0(_173_),
    .S1(_174_),
    .X(_176_));
 sky130_fd_sc_hd__clkbuf_1 _450_ (.A(_176_),
    .X(net53));
 sky130_fd_sc_hd__mux4_1 _451_ (.A0(\memblk.FIFO[0][25] ),
    .A1(\memblk.FIFO[1][25] ),
    .A2(\memblk.FIFO[2][25] ),
    .A3(\memblk.FIFO[3][25] ),
    .S0(_173_),
    .S1(_174_),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_1 _452_ (.A(_177_),
    .X(net54));
 sky130_fd_sc_hd__mux4_1 _453_ (.A0(\memblk.FIFO[0][26] ),
    .A1(\memblk.FIFO[1][26] ),
    .A2(\memblk.FIFO[2][26] ),
    .A3(\memblk.FIFO[3][26] ),
    .S0(_173_),
    .S1(_174_),
    .X(_178_));
 sky130_fd_sc_hd__clkbuf_1 _454_ (.A(_178_),
    .X(net55));
 sky130_fd_sc_hd__mux4_1 _455_ (.A0(\memblk.FIFO[0][27] ),
    .A1(\memblk.FIFO[1][27] ),
    .A2(\memblk.FIFO[2][27] ),
    .A3(\memblk.FIFO[3][27] ),
    .S0(_173_),
    .S1(_174_),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_1 _456_ (.A(_179_),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 _457_ (.A0(\memblk.FIFO[0][28] ),
    .A1(\memblk.FIFO[1][28] ),
    .A2(\memblk.FIFO[2][28] ),
    .A3(\memblk.FIFO[3][28] ),
    .S0(_173_),
    .S1(_174_),
    .X(_180_));
 sky130_fd_sc_hd__clkbuf_1 _458_ (.A(_180_),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 _459_ (.A0(\memblk.FIFO[0][29] ),
    .A1(\memblk.FIFO[1][29] ),
    .A2(\memblk.FIFO[2][29] ),
    .A3(\memblk.FIFO[3][29] ),
    .S0(_140_),
    .S1(_142_),
    .X(_181_));
 sky130_fd_sc_hd__clkbuf_1 _460_ (.A(_181_),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 _461_ (.A0(\memblk.FIFO[0][30] ),
    .A1(\memblk.FIFO[1][30] ),
    .A2(\memblk.FIFO[2][30] ),
    .A3(\memblk.FIFO[3][30] ),
    .S0(_140_),
    .S1(_142_),
    .X(_182_));
 sky130_fd_sc_hd__clkbuf_1 _462_ (.A(_182_),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 _463_ (.A0(\memblk.FIFO[0][31] ),
    .A1(\memblk.FIFO[1][31] ),
    .A2(\memblk.FIFO[2][31] ),
    .A3(\memblk.FIFO[3][31] ),
    .S0(_140_),
    .S1(_142_),
    .X(_183_));
 sky130_fd_sc_hd__clkbuf_1 _464_ (.A(_183_),
    .X(net61));
 sky130_fd_sc_hd__or3b_1 _465_ (.A(net34),
    .B(\memblk.wr_addr[0] ),
    .C_N(\memblk.wr_addr[1] ),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_2 _466_ (.A(_184_),
    .X(_185_));
 sky130_fd_sc_hd__buf_2 _467_ (.A(_185_),
    .X(_186_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(net1),
    .A1(net112),
    .S(_186_),
    .X(_187_));
 sky130_fd_sc_hd__clkbuf_1 _469_ (.A(_187_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(net12),
    .A1(net191),
    .S(_186_),
    .X(_188_));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(_188_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(net23),
    .A1(net186),
    .S(_186_),
    .X(_189_));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(_189_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(net26),
    .A1(net122),
    .S(_186_),
    .X(_190_));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(_190_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(net27),
    .A1(net124),
    .S(_186_),
    .X(_191_));
 sky130_fd_sc_hd__clkbuf_1 _477_ (.A(_191_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _478_ (.A0(net28),
    .A1(net134),
    .S(_186_),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(_192_),
    .X(_005_));
 sky130_fd_sc_hd__buf_2 _480_ (.A(_185_),
    .X(_193_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(net29),
    .A1(net139),
    .S(_193_),
    .X(_194_));
 sky130_fd_sc_hd__clkbuf_1 _482_ (.A(_194_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(net30),
    .A1(net187),
    .S(_193_),
    .X(_195_));
 sky130_fd_sc_hd__clkbuf_1 _484_ (.A(_195_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(net31),
    .A1(net183),
    .S(_193_),
    .X(_196_));
 sky130_fd_sc_hd__clkbuf_1 _486_ (.A(_196_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(net32),
    .A1(net103),
    .S(_193_),
    .X(_197_));
 sky130_fd_sc_hd__clkbuf_1 _488_ (.A(_197_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _489_ (.A0(net2),
    .A1(net114),
    .S(_193_),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _490_ (.A(_198_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(net3),
    .A1(net107),
    .S(_193_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_1 _492_ (.A(_199_),
    .X(_011_));
 sky130_fd_sc_hd__buf_2 _493_ (.A(_185_),
    .X(_200_));
 sky130_fd_sc_hd__mux2_1 _494_ (.A0(net4),
    .A1(net95),
    .S(_200_),
    .X(_201_));
 sky130_fd_sc_hd__clkbuf_1 _495_ (.A(_201_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _496_ (.A0(net5),
    .A1(net125),
    .S(_200_),
    .X(_202_));
 sky130_fd_sc_hd__clkbuf_1 _497_ (.A(_202_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _498_ (.A0(net6),
    .A1(net102),
    .S(_200_),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(_203_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _500_ (.A0(net7),
    .A1(net167),
    .S(_200_),
    .X(_204_));
 sky130_fd_sc_hd__clkbuf_1 _501_ (.A(_204_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _502_ (.A0(net8),
    .A1(net171),
    .S(_200_),
    .X(_205_));
 sky130_fd_sc_hd__clkbuf_1 _503_ (.A(_205_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _504_ (.A0(net9),
    .A1(net185),
    .S(_200_),
    .X(_206_));
 sky130_fd_sc_hd__clkbuf_1 _505_ (.A(_206_),
    .X(_017_));
 sky130_fd_sc_hd__buf_2 _506_ (.A(_185_),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _507_ (.A0(net10),
    .A1(net174),
    .S(_207_),
    .X(_208_));
 sky130_fd_sc_hd__clkbuf_1 _508_ (.A(_208_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _509_ (.A0(net11),
    .A1(net190),
    .S(_207_),
    .X(_209_));
 sky130_fd_sc_hd__clkbuf_1 _510_ (.A(_209_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _511_ (.A0(net13),
    .A1(net123),
    .S(_207_),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_1 _512_ (.A(_210_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _513_ (.A0(net14),
    .A1(net164),
    .S(_207_),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _514_ (.A(_211_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _515_ (.A0(net15),
    .A1(net157),
    .S(_207_),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_1 _516_ (.A(_212_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _517_ (.A0(net16),
    .A1(net113),
    .S(_207_),
    .X(_213_));
 sky130_fd_sc_hd__clkbuf_1 _518_ (.A(_213_),
    .X(_023_));
 sky130_fd_sc_hd__buf_2 _519_ (.A(_184_),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _520_ (.A0(net17),
    .A1(net117),
    .S(_214_),
    .X(_215_));
 sky130_fd_sc_hd__clkbuf_1 _521_ (.A(_215_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _522_ (.A0(net18),
    .A1(net146),
    .S(_214_),
    .X(_216_));
 sky130_fd_sc_hd__clkbuf_1 _523_ (.A(_216_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _524_ (.A0(net19),
    .A1(net179),
    .S(_214_),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_1 _525_ (.A(_217_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _526_ (.A0(net20),
    .A1(net155),
    .S(_214_),
    .X(_218_));
 sky130_fd_sc_hd__clkbuf_1 _527_ (.A(_218_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _528_ (.A0(net21),
    .A1(net198),
    .S(_214_),
    .X(_219_));
 sky130_fd_sc_hd__clkbuf_1 _529_ (.A(_219_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _530_ (.A0(net22),
    .A1(net147),
    .S(_214_),
    .X(_220_));
 sky130_fd_sc_hd__clkbuf_1 _531_ (.A(_220_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _532_ (.A0(net24),
    .A1(net142),
    .S(_185_),
    .X(_221_));
 sky130_fd_sc_hd__clkbuf_1 _533_ (.A(_221_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _534_ (.A0(net25),
    .A1(net188),
    .S(_185_),
    .X(_222_));
 sky130_fd_sc_hd__clkbuf_1 _535_ (.A(_222_),
    .X(_031_));
 sky130_fd_sc_hd__clkbuf_2 _536_ (.A(net33),
    .X(_223_));
 sky130_fd_sc_hd__nand2b_1 _537_ (.A_N(net34),
    .B(\memblk.wr_addr[0] ),
    .Y(_224_));
 sky130_fd_sc_hd__inv_1 _538_ (.A(net34),
    .Y(_225_));
 sky130_fd_sc_hd__or2_1 _539_ (.A(_225_),
    .B(\memblk.wr_addr[0] ),
    .X(_226_));
 sky130_fd_sc_hd__and3_1 _540_ (.A(_223_),
    .B(_224_),
    .C(_226_),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(_227_),
    .X(_032_));
 sky130_fd_sc_hd__or2_1 _542_ (.A(\memblk.wr_addr[1] ),
    .B(_224_),
    .X(_228_));
 sky130_fd_sc_hd__clkbuf_2 _543_ (.A(_228_),
    .X(_229_));
 sky130_fd_sc_hd__buf_2 _544_ (.A(_229_),
    .X(_230_));
 sky130_fd_sc_hd__nand2_1 _545_ (.A(net204),
    .B(_224_),
    .Y(_231_));
 sky130_fd_sc_hd__inv_2 _546_ (.A(_223_),
    .Y(_232_));
 sky130_fd_sc_hd__a21oi_1 _547_ (.A1(_230_),
    .A2(_231_),
    .B1(_232_),
    .Y(_033_));
 sky130_fd_sc_hd__or3_1 _548_ (.A(net34),
    .B(\memblk.wr_addr[0] ),
    .C(\memblk.wr_addr[1] ),
    .X(_233_));
 sky130_fd_sc_hd__clkbuf_2 _549_ (.A(_233_),
    .X(_234_));
 sky130_fd_sc_hd__buf_2 _550_ (.A(_234_),
    .X(_235_));
 sky130_fd_sc_hd__mux2_1 _551_ (.A0(net1),
    .A1(net176),
    .S(_235_),
    .X(_236_));
 sky130_fd_sc_hd__clkbuf_1 _552_ (.A(_236_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(net12),
    .A1(net133),
    .S(_235_),
    .X(_237_));
 sky130_fd_sc_hd__clkbuf_1 _554_ (.A(_237_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(net23),
    .A1(net129),
    .S(_235_),
    .X(_238_));
 sky130_fd_sc_hd__clkbuf_1 _556_ (.A(_238_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _557_ (.A0(net26),
    .A1(net199),
    .S(_235_),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _558_ (.A(_239_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _559_ (.A0(net27),
    .A1(net144),
    .S(_235_),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_1 _560_ (.A(_240_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _561_ (.A0(net28),
    .A1(net178),
    .S(_235_),
    .X(_241_));
 sky130_fd_sc_hd__clkbuf_1 _562_ (.A(_241_),
    .X(_039_));
 sky130_fd_sc_hd__buf_2 _563_ (.A(_234_),
    .X(_242_));
 sky130_fd_sc_hd__mux2_1 _564_ (.A0(net29),
    .A1(net156),
    .S(_242_),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _565_ (.A(_243_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _566_ (.A0(net30),
    .A1(net121),
    .S(_242_),
    .X(_244_));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(_244_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _568_ (.A0(net31),
    .A1(net115),
    .S(_242_),
    .X(_245_));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(_245_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _570_ (.A0(net32),
    .A1(net87),
    .S(_242_),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(_246_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _572_ (.A0(net2),
    .A1(net106),
    .S(_242_),
    .X(_247_));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(_247_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _574_ (.A0(net3),
    .A1(net170),
    .S(_242_),
    .X(_248_));
 sky130_fd_sc_hd__clkbuf_1 _575_ (.A(_248_),
    .X(_045_));
 sky130_fd_sc_hd__buf_2 _576_ (.A(_234_),
    .X(_249_));
 sky130_fd_sc_hd__mux2_1 _577_ (.A0(net4),
    .A1(net111),
    .S(_249_),
    .X(_250_));
 sky130_fd_sc_hd__clkbuf_1 _578_ (.A(_250_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _579_ (.A0(net5),
    .A1(net194),
    .S(_249_),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_1 _580_ (.A(_251_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _581_ (.A0(net6),
    .A1(net193),
    .S(_249_),
    .X(_252_));
 sky130_fd_sc_hd__clkbuf_1 _582_ (.A(_252_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _583_ (.A0(net7),
    .A1(net138),
    .S(_249_),
    .X(_253_));
 sky130_fd_sc_hd__clkbuf_1 _584_ (.A(_253_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _585_ (.A0(net8),
    .A1(net180),
    .S(_249_),
    .X(_254_));
 sky130_fd_sc_hd__clkbuf_1 _586_ (.A(_254_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _587_ (.A0(net9),
    .A1(net158),
    .S(_249_),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _588_ (.A(_255_),
    .X(_051_));
 sky130_fd_sc_hd__buf_2 _589_ (.A(_234_),
    .X(_256_));
 sky130_fd_sc_hd__mux2_1 _590_ (.A0(net10),
    .A1(net201),
    .S(_256_),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _591_ (.A(_257_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _592_ (.A0(net11),
    .A1(net160),
    .S(_256_),
    .X(_258_));
 sky130_fd_sc_hd__clkbuf_1 _593_ (.A(_258_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _594_ (.A0(net13),
    .A1(net168),
    .S(_256_),
    .X(_259_));
 sky130_fd_sc_hd__clkbuf_1 _595_ (.A(_259_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _596_ (.A0(net14),
    .A1(net141),
    .S(_256_),
    .X(_260_));
 sky130_fd_sc_hd__clkbuf_1 _597_ (.A(_260_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _598_ (.A0(net15),
    .A1(net150),
    .S(_256_),
    .X(_261_));
 sky130_fd_sc_hd__clkbuf_1 _599_ (.A(_261_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _600_ (.A0(net16),
    .A1(net105),
    .S(_256_),
    .X(_262_));
 sky130_fd_sc_hd__clkbuf_1 _601_ (.A(_262_),
    .X(_057_));
 sky130_fd_sc_hd__buf_2 _602_ (.A(_233_),
    .X(_263_));
 sky130_fd_sc_hd__mux2_1 _603_ (.A0(net17),
    .A1(net137),
    .S(_263_),
    .X(_264_));
 sky130_fd_sc_hd__clkbuf_1 _604_ (.A(_264_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _605_ (.A0(net18),
    .A1(net189),
    .S(_263_),
    .X(_265_));
 sky130_fd_sc_hd__clkbuf_1 _606_ (.A(_265_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _607_ (.A0(net19),
    .A1(net166),
    .S(_263_),
    .X(_266_));
 sky130_fd_sc_hd__clkbuf_1 _608_ (.A(_266_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _609_ (.A0(net20),
    .A1(net120),
    .S(_263_),
    .X(_267_));
 sky130_fd_sc_hd__clkbuf_1 _610_ (.A(_267_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _611_ (.A0(net21),
    .A1(net203),
    .S(_263_),
    .X(_268_));
 sky130_fd_sc_hd__clkbuf_1 _612_ (.A(_268_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _613_ (.A0(net22),
    .A1(net192),
    .S(_263_),
    .X(_269_));
 sky130_fd_sc_hd__clkbuf_1 _614_ (.A(_269_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _615_ (.A0(net24),
    .A1(net163),
    .S(_234_),
    .X(_270_));
 sky130_fd_sc_hd__clkbuf_1 _616_ (.A(_270_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _617_ (.A0(net25),
    .A1(net169),
    .S(_234_),
    .X(_271_));
 sky130_fd_sc_hd__clkbuf_1 _618_ (.A(_271_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _619_ (.A0(net1),
    .A1(net90),
    .S(_230_),
    .X(_272_));
 sky130_fd_sc_hd__clkbuf_1 _620_ (.A(_272_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _621_ (.A0(net12),
    .A1(net177),
    .S(_230_),
    .X(_273_));
 sky130_fd_sc_hd__clkbuf_1 _622_ (.A(_273_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _623_ (.A0(net23),
    .A1(net148),
    .S(_230_),
    .X(_274_));
 sky130_fd_sc_hd__clkbuf_1 _624_ (.A(_274_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _625_ (.A0(net26),
    .A1(net195),
    .S(_230_),
    .X(_275_));
 sky130_fd_sc_hd__clkbuf_1 _626_ (.A(_275_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _627_ (.A0(net27),
    .A1(net110),
    .S(_230_),
    .X(_276_));
 sky130_fd_sc_hd__clkbuf_1 _628_ (.A(_276_),
    .X(_070_));
 sky130_fd_sc_hd__buf_2 _629_ (.A(_229_),
    .X(_277_));
 sky130_fd_sc_hd__mux2_1 _630_ (.A0(net28),
    .A1(net165),
    .S(_277_),
    .X(_278_));
 sky130_fd_sc_hd__clkbuf_1 _631_ (.A(_278_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _632_ (.A0(net29),
    .A1(net149),
    .S(_277_),
    .X(_279_));
 sky130_fd_sc_hd__clkbuf_1 _633_ (.A(_279_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _634_ (.A0(net30),
    .A1(net153),
    .S(_277_),
    .X(_280_));
 sky130_fd_sc_hd__clkbuf_1 _635_ (.A(_280_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _636_ (.A0(net31),
    .A1(net162),
    .S(_277_),
    .X(_281_));
 sky130_fd_sc_hd__clkbuf_1 _637_ (.A(_281_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _638_ (.A0(net32),
    .A1(net132),
    .S(_277_),
    .X(_282_));
 sky130_fd_sc_hd__clkbuf_1 _639_ (.A(_282_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _640_ (.A0(net2),
    .A1(net104),
    .S(_277_),
    .X(_283_));
 sky130_fd_sc_hd__clkbuf_1 _641_ (.A(_283_),
    .X(_076_));
 sky130_fd_sc_hd__buf_2 _642_ (.A(_229_),
    .X(_284_));
 sky130_fd_sc_hd__mux2_1 _643_ (.A0(net3),
    .A1(net173),
    .S(_284_),
    .X(_285_));
 sky130_fd_sc_hd__clkbuf_1 _644_ (.A(_285_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _645_ (.A0(net4),
    .A1(net143),
    .S(_284_),
    .X(_286_));
 sky130_fd_sc_hd__clkbuf_1 _646_ (.A(_286_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _647_ (.A0(net5),
    .A1(net161),
    .S(_284_),
    .X(_287_));
 sky130_fd_sc_hd__clkbuf_1 _648_ (.A(_287_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _649_ (.A0(net6),
    .A1(net126),
    .S(_284_),
    .X(_288_));
 sky130_fd_sc_hd__clkbuf_1 _650_ (.A(_288_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _651_ (.A0(net7),
    .A1(net175),
    .S(_284_),
    .X(_289_));
 sky130_fd_sc_hd__clkbuf_1 _652_ (.A(_289_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _653_ (.A0(net8),
    .A1(net196),
    .S(_284_),
    .X(_290_));
 sky130_fd_sc_hd__clkbuf_1 _654_ (.A(_290_),
    .X(_082_));
 sky130_fd_sc_hd__buf_2 _655_ (.A(_228_),
    .X(_291_));
 sky130_fd_sc_hd__mux2_1 _656_ (.A0(net9),
    .A1(net152),
    .S(_291_),
    .X(_292_));
 sky130_fd_sc_hd__clkbuf_1 _657_ (.A(_292_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _658_ (.A0(net10),
    .A1(net136),
    .S(_291_),
    .X(_293_));
 sky130_fd_sc_hd__clkbuf_1 _659_ (.A(_293_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _660_ (.A0(net11),
    .A1(net151),
    .S(_291_),
    .X(_294_));
 sky130_fd_sc_hd__clkbuf_1 _661_ (.A(_294_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _662_ (.A0(net13),
    .A1(net172),
    .S(_291_),
    .X(_295_));
 sky130_fd_sc_hd__clkbuf_1 _663_ (.A(_295_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _664_ (.A0(net14),
    .A1(net93),
    .S(_291_),
    .X(_296_));
 sky130_fd_sc_hd__clkbuf_1 _665_ (.A(_296_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _666_ (.A0(net15),
    .A1(net140),
    .S(_291_),
    .X(_297_));
 sky130_fd_sc_hd__clkbuf_1 _667_ (.A(_297_),
    .X(_088_));
 sky130_fd_sc_hd__buf_2 _668_ (.A(_228_),
    .X(_298_));
 sky130_fd_sc_hd__mux2_1 _669_ (.A0(net16),
    .A1(net91),
    .S(_298_),
    .X(_299_));
 sky130_fd_sc_hd__clkbuf_1 _670_ (.A(_299_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _671_ (.A0(net17),
    .A1(net135),
    .S(_298_),
    .X(_300_));
 sky130_fd_sc_hd__clkbuf_1 _672_ (.A(_300_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _673_ (.A0(net18),
    .A1(net200),
    .S(_298_),
    .X(_301_));
 sky130_fd_sc_hd__clkbuf_1 _674_ (.A(_301_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _675_ (.A0(net19),
    .A1(net159),
    .S(_298_),
    .X(_302_));
 sky130_fd_sc_hd__clkbuf_1 _676_ (.A(_302_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _677_ (.A0(net20),
    .A1(net181),
    .S(_298_),
    .X(_303_));
 sky130_fd_sc_hd__clkbuf_1 _678_ (.A(_303_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _679_ (.A0(net21),
    .A1(net154),
    .S(_298_),
    .X(_304_));
 sky130_fd_sc_hd__clkbuf_1 _680_ (.A(_304_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _681_ (.A0(net22),
    .A1(net182),
    .S(_229_),
    .X(_305_));
 sky130_fd_sc_hd__clkbuf_1 _682_ (.A(_305_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _683_ (.A0(net24),
    .A1(net197),
    .S(_229_),
    .X(_306_));
 sky130_fd_sc_hd__clkbuf_1 _684_ (.A(_306_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _685_ (.A0(net25),
    .A1(net202),
    .S(_229_),
    .X(_307_));
 sky130_fd_sc_hd__clkbuf_1 _686_ (.A(_307_),
    .X(_097_));
 sky130_fd_sc_hd__and3_1 _687_ (.A(_225_),
    .B(\memblk.wr_addr[0] ),
    .C(\memblk.wr_addr[1] ),
    .X(_308_));
 sky130_fd_sc_hd__clkbuf_2 _688_ (.A(_308_),
    .X(_309_));
 sky130_fd_sc_hd__buf_2 _689_ (.A(_309_),
    .X(_310_));
 sky130_fd_sc_hd__mux2_1 _690_ (.A0(net86),
    .A1(net1),
    .S(_310_),
    .X(_311_));
 sky130_fd_sc_hd__clkbuf_1 _691_ (.A(_311_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _692_ (.A0(net128),
    .A1(net12),
    .S(_310_),
    .X(_312_));
 sky130_fd_sc_hd__clkbuf_1 _693_ (.A(_312_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _694_ (.A0(net82),
    .A1(net23),
    .S(_310_),
    .X(_313_));
 sky130_fd_sc_hd__clkbuf_1 _695_ (.A(_313_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _696_ (.A0(net80),
    .A1(net26),
    .S(_310_),
    .X(_314_));
 sky130_fd_sc_hd__clkbuf_1 _697_ (.A(_314_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _698_ (.A0(net83),
    .A1(net27),
    .S(_310_),
    .X(_315_));
 sky130_fd_sc_hd__clkbuf_1 _699_ (.A(_315_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _700_ (.A0(net131),
    .A1(net28),
    .S(_310_),
    .X(_316_));
 sky130_fd_sc_hd__clkbuf_1 _701_ (.A(_316_),
    .X(_103_));
 sky130_fd_sc_hd__buf_2 _702_ (.A(_309_),
    .X(_317_));
 sky130_fd_sc_hd__mux2_1 _703_ (.A0(net97),
    .A1(net29),
    .S(_317_),
    .X(_318_));
 sky130_fd_sc_hd__clkbuf_1 _704_ (.A(_318_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _705_ (.A0(net78),
    .A1(net30),
    .S(_317_),
    .X(_319_));
 sky130_fd_sc_hd__clkbuf_1 _706_ (.A(_319_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _707_ (.A0(net85),
    .A1(net31),
    .S(_317_),
    .X(_320_));
 sky130_fd_sc_hd__clkbuf_1 _708_ (.A(_320_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _709_ (.A0(net101),
    .A1(net32),
    .S(_317_),
    .X(_321_));
 sky130_fd_sc_hd__clkbuf_1 _710_ (.A(_321_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _711_ (.A0(net96),
    .A1(net2),
    .S(_317_),
    .X(_322_));
 sky130_fd_sc_hd__clkbuf_1 _712_ (.A(_322_),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _713_ (.A0(net118),
    .A1(net3),
    .S(_317_),
    .X(_323_));
 sky130_fd_sc_hd__clkbuf_1 _714_ (.A(_323_),
    .X(_109_));
 sky130_fd_sc_hd__buf_2 _715_ (.A(_309_),
    .X(_324_));
 sky130_fd_sc_hd__mux2_1 _716_ (.A0(net145),
    .A1(net4),
    .S(_324_),
    .X(_325_));
 sky130_fd_sc_hd__clkbuf_1 _717_ (.A(_325_),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _718_ (.A0(net88),
    .A1(net5),
    .S(_324_),
    .X(_326_));
 sky130_fd_sc_hd__clkbuf_1 _719_ (.A(_326_),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _720_ (.A0(net130),
    .A1(net6),
    .S(_324_),
    .X(_327_));
 sky130_fd_sc_hd__clkbuf_1 _721_ (.A(_327_),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _722_ (.A0(net76),
    .A1(net7),
    .S(_324_),
    .X(_328_));
 sky130_fd_sc_hd__clkbuf_1 _723_ (.A(_328_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _724_ (.A0(net116),
    .A1(net8),
    .S(_324_),
    .X(_329_));
 sky130_fd_sc_hd__clkbuf_1 _725_ (.A(_329_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _726_ (.A0(net98),
    .A1(net9),
    .S(_324_),
    .X(_330_));
 sky130_fd_sc_hd__clkbuf_1 _727_ (.A(_330_),
    .X(_115_));
 sky130_fd_sc_hd__buf_2 _728_ (.A(_309_),
    .X(_331_));
 sky130_fd_sc_hd__mux2_1 _729_ (.A0(net81),
    .A1(net10),
    .S(_331_),
    .X(_332_));
 sky130_fd_sc_hd__clkbuf_1 _730_ (.A(_332_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _731_ (.A0(net92),
    .A1(net11),
    .S(_331_),
    .X(_333_));
 sky130_fd_sc_hd__clkbuf_1 _732_ (.A(_333_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _733_ (.A0(net84),
    .A1(net13),
    .S(_331_),
    .X(_334_));
 sky130_fd_sc_hd__clkbuf_1 _734_ (.A(_334_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _735_ (.A0(net184),
    .A1(net14),
    .S(_331_),
    .X(_335_));
 sky130_fd_sc_hd__clkbuf_1 _736_ (.A(_335_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _737_ (.A0(net119),
    .A1(net15),
    .S(_331_),
    .X(_336_));
 sky130_fd_sc_hd__clkbuf_1 _738_ (.A(_336_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _739_ (.A0(net100),
    .A1(net16),
    .S(_331_),
    .X(_337_));
 sky130_fd_sc_hd__clkbuf_1 _740_ (.A(_337_),
    .X(_121_));
 sky130_fd_sc_hd__buf_2 _741_ (.A(_308_),
    .X(_338_));
 sky130_fd_sc_hd__mux2_1 _742_ (.A0(net108),
    .A1(net17),
    .S(_338_),
    .X(_339_));
 sky130_fd_sc_hd__clkbuf_1 _743_ (.A(_339_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _744_ (.A0(net89),
    .A1(net18),
    .S(_338_),
    .X(_340_));
 sky130_fd_sc_hd__clkbuf_1 _745_ (.A(_340_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _746_ (.A0(net127),
    .A1(net19),
    .S(_338_),
    .X(_341_));
 sky130_fd_sc_hd__clkbuf_1 _747_ (.A(_341_),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _748_ (.A0(net77),
    .A1(net20),
    .S(_338_),
    .X(_342_));
 sky130_fd_sc_hd__clkbuf_1 _749_ (.A(_342_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _750_ (.A0(net99),
    .A1(net21),
    .S(_338_),
    .X(_343_));
 sky130_fd_sc_hd__clkbuf_1 _751_ (.A(_343_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _752_ (.A0(net109),
    .A1(net22),
    .S(_338_),
    .X(_344_));
 sky130_fd_sc_hd__clkbuf_1 _753_ (.A(_344_),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _754_ (.A0(net94),
    .A1(net24),
    .S(_309_),
    .X(_345_));
 sky130_fd_sc_hd__clkbuf_1 _755_ (.A(_345_),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _756_ (.A0(net79),
    .A1(net25),
    .S(_309_),
    .X(_346_));
 sky130_fd_sc_hd__clkbuf_1 _757_ (.A(_346_),
    .X(_129_));
 sky130_fd_sc_hd__inv_2 _758_ (.A(net35),
    .Y(_347_));
 sky130_fd_sc_hd__buf_6 _759_ (.A(net34),
    .X(_348_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _760_ (.A(_348_),
    .X(_349_));
 sky130_fd_sc_hd__o21ai_1 _761_ (.A1(net72),
    .A2(_349_),
    .B1(net71),
    .Y(_350_));
 sky130_fd_sc_hd__or3b_1 _762_ (.A(_347_),
    .B(_232_),
    .C_N(_350_),
    .X(_351_));
 sky130_fd_sc_hd__clkbuf_1 _763_ (.A(_351_),
    .X(_130_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _764_ (.A(net35),
    .X(_352_));
 sky130_fd_sc_hd__nor2_1 _765_ (.A(_352_),
    .B(_350_),
    .Y(_353_));
 sky130_fd_sc_hd__buf_1 _766_ (.A(\fcounter[0] ),
    .X(_354_));
 sky130_fd_sc_hd__or4b_1 _767_ (.A(_348_),
    .B(_354_),
    .C(\fcounter[2] ),
    .D_N(\fcounter[1] ),
    .X(_355_));
 sky130_fd_sc_hd__o211a_1 _768_ (.A1(net72),
    .A2(_225_),
    .B1(_355_),
    .C1(_352_),
    .X(_356_));
 sky130_fd_sc_hd__or3_1 _769_ (.A(_232_),
    .B(_353_),
    .C(_356_),
    .X(_357_));
 sky130_fd_sc_hd__clkbuf_1 _770_ (.A(_357_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _771_ (.A0(net73),
    .A1(net72),
    .S(_349_),
    .X(_358_));
 sky130_fd_sc_hd__buf_1 _772_ (.A(\fcounter[2] ),
    .X(_359_));
 sky130_fd_sc_hd__or4b_1 _773_ (.A(_348_),
    .B(\fcounter[1] ),
    .C(_359_),
    .D_N(_354_),
    .X(_360_));
 sky130_fd_sc_hd__o211a_1 _774_ (.A1(_225_),
    .A2(net73),
    .B1(_360_),
    .C1(_352_),
    .X(_361_));
 sky130_fd_sc_hd__a211o_1 _775_ (.A1(_347_),
    .A2(_358_),
    .B1(_361_),
    .C1(_232_),
    .X(_132_));
 sky130_fd_sc_hd__inv_2 _776_ (.A(net70),
    .Y(_362_));
 sky130_fd_sc_hd__nor2_1 _777_ (.A(_349_),
    .B(net69),
    .Y(_363_));
 sky130_fd_sc_hd__a31o_1 _778_ (.A1(_352_),
    .A2(_349_),
    .A3(_362_),
    .B1(_363_),
    .X(_364_));
 sky130_fd_sc_hd__nand4bb_1 _779_ (.A_N(_354_),
    .B_N(_359_),
    .C(_349_),
    .D(\fcounter[1] ),
    .Y(_365_));
 sky130_fd_sc_hd__or2_1 _780_ (.A(_349_),
    .B(net70),
    .X(_366_));
 sky130_fd_sc_hd__a21oi_1 _781_ (.A1(_365_),
    .A2(_366_),
    .B1(_352_),
    .Y(_367_));
 sky130_fd_sc_hd__o21ai_1 _782_ (.A1(_364_),
    .A2(_367_),
    .B1(_223_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2_1 _783_ (.A0(net69),
    .A1(_363_),
    .S(_223_),
    .X(_368_));
 sky130_fd_sc_hd__clkbuf_1 _784_ (.A(_368_),
    .X(_134_));
 sky130_fd_sc_hd__and2_1 _785_ (.A(_223_),
    .B(_354_),
    .X(_369_));
 sky130_fd_sc_hd__nor2_1 _786_ (.A(_232_),
    .B(_354_),
    .Y(_370_));
 sky130_fd_sc_hd__and3b_1 _787_ (.A_N(net35),
    .B(_348_),
    .C(net69),
    .X(_371_));
 sky130_fd_sc_hd__a31o_1 _788_ (.A1(net71),
    .A2(net35),
    .A3(_225_),
    .B1(_371_),
    .X(_372_));
 sky130_fd_sc_hd__mux2_1 _789_ (.A0(_369_),
    .A1(_370_),
    .S(_372_),
    .X(_373_));
 sky130_fd_sc_hd__clkbuf_1 _790_ (.A(_373_),
    .X(_135_));
 sky130_fd_sc_hd__and2b_1 _791_ (.A_N(\fcounter[1] ),
    .B(net33),
    .X(_374_));
 sky130_fd_sc_hd__and2_1 _792_ (.A(net33),
    .B(\fcounter[1] ),
    .X(_375_));
 sky130_fd_sc_hd__and4bb_1 _793_ (.A_N(net35),
    .B_N(\fcounter[0] ),
    .C(net69),
    .D(_348_),
    .X(_376_));
 sky130_fd_sc_hd__and4b_1 _794_ (.A_N(_348_),
    .B(_354_),
    .C(net71),
    .D(net35),
    .X(_377_));
 sky130_fd_sc_hd__nor2_1 _795_ (.A(_376_),
    .B(_377_),
    .Y(_378_));
 sky130_fd_sc_hd__mux2_1 _796_ (.A0(_374_),
    .A1(_375_),
    .S(_378_),
    .X(_379_));
 sky130_fd_sc_hd__clkbuf_1 _797_ (.A(_379_),
    .X(_136_));
 sky130_fd_sc_hd__and3b_1 _798_ (.A_N(_377_),
    .B(_375_),
    .C(_359_),
    .X(_380_));
 sky130_fd_sc_hd__and3b_1 _799_ (.A_N(_359_),
    .B(_377_),
    .C(_375_),
    .X(_381_));
 sky130_fd_sc_hd__and3b_1 _800_ (.A_N(_376_),
    .B(_374_),
    .C(_359_),
    .X(_382_));
 sky130_fd_sc_hd__and3b_1 _801_ (.A_N(_359_),
    .B(_376_),
    .C(_374_),
    .X(_383_));
 sky130_fd_sc_hd__or4_1 _802_ (.A(_380_),
    .B(_381_),
    .C(_382_),
    .D(_383_),
    .X(_384_));
 sky130_fd_sc_hd__clkbuf_1 _803_ (.A(_384_),
    .X(_137_));
 sky130_fd_sc_hd__or2b_1 _804_ (.A(_352_),
    .B_N(_140_),
    .X(_385_));
 sky130_fd_sc_hd__or2_1 _805_ (.A(_347_),
    .B(_141_),
    .X(_386_));
 sky130_fd_sc_hd__and3_1 _806_ (.A(_223_),
    .B(_385_),
    .C(_386_),
    .X(_387_));
 sky130_fd_sc_hd__clkbuf_1 _807_ (.A(_387_),
    .X(_138_));
 sky130_fd_sc_hd__xor2_1 _808_ (.A(_143_),
    .B(_385_),
    .X(_388_));
 sky130_fd_sc_hd__nor2_1 _809_ (.A(_232_),
    .B(_388_),
    .Y(_139_));
 sky130_fd_sc_hd__dfxtp_1 _810_ (.CLK(clknet_4_1_0_Clk),
    .D(_000_),
    .Q(\memblk.FIFO[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _811_ (.CLK(clknet_4_0_0_Clk),
    .D(_001_),
    .Q(\memblk.FIFO[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _812_ (.CLK(clknet_4_0_0_Clk),
    .D(_002_),
    .Q(\memblk.FIFO[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _813_ (.CLK(clknet_4_0_0_Clk),
    .D(_003_),
    .Q(\memblk.FIFO[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _814_ (.CLK(clknet_4_3_0_Clk),
    .D(_004_),
    .Q(\memblk.FIFO[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _815_ (.CLK(clknet_4_1_0_Clk),
    .D(_005_),
    .Q(\memblk.FIFO[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _816_ (.CLK(clknet_4_4_0_Clk),
    .D(_006_),
    .Q(\memblk.FIFO[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _817_ (.CLK(clknet_4_5_0_Clk),
    .D(_007_),
    .Q(\memblk.FIFO[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _818_ (.CLK(clknet_4_4_0_Clk),
    .D(_008_),
    .Q(\memblk.FIFO[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _819_ (.CLK(clknet_4_4_0_Clk),
    .D(_009_),
    .Q(\memblk.FIFO[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _820_ (.CLK(clknet_4_4_0_Clk),
    .D(_010_),
    .Q(\memblk.FIFO[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _821_ (.CLK(clknet_4_5_0_Clk),
    .D(_011_),
    .Q(\memblk.FIFO[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _822_ (.CLK(clknet_4_6_0_Clk),
    .D(_012_),
    .Q(\memblk.FIFO[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _823_ (.CLK(clknet_4_7_0_Clk),
    .D(_013_),
    .Q(\memblk.FIFO[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _824_ (.CLK(clknet_4_13_0_Clk),
    .D(_014_),
    .Q(\memblk.FIFO[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _825_ (.CLK(clknet_4_7_0_Clk),
    .D(_015_),
    .Q(\memblk.FIFO[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _826_ (.CLK(clknet_4_13_0_Clk),
    .D(_016_),
    .Q(\memblk.FIFO[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _827_ (.CLK(clknet_4_12_0_Clk),
    .D(_017_),
    .Q(\memblk.FIFO[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _828_ (.CLK(clknet_4_9_0_Clk),
    .D(_018_),
    .Q(\memblk.FIFO[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _829_ (.CLK(clknet_4_14_0_Clk),
    .D(_019_),
    .Q(\memblk.FIFO[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _830_ (.CLK(clknet_4_14_0_Clk),
    .D(_020_),
    .Q(\memblk.FIFO[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _831_ (.CLK(clknet_4_15_0_Clk),
    .D(_021_),
    .Q(\memblk.FIFO[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _832_ (.CLK(clknet_4_12_0_Clk),
    .D(_022_),
    .Q(\memblk.FIFO[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _833_ (.CLK(clknet_4_11_0_Clk),
    .D(_023_),
    .Q(\memblk.FIFO[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _834_ (.CLK(clknet_4_9_0_Clk),
    .D(_024_),
    .Q(\memblk.FIFO[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _835_ (.CLK(clknet_4_8_0_Clk),
    .D(_025_),
    .Q(\memblk.FIFO[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _836_ (.CLK(clknet_4_10_0_Clk),
    .D(_026_),
    .Q(\memblk.FIFO[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _837_ (.CLK(clknet_4_8_0_Clk),
    .D(_027_),
    .Q(\memblk.FIFO[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _838_ (.CLK(clknet_4_10_0_Clk),
    .D(_028_),
    .Q(\memblk.FIFO[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _839_ (.CLK(clknet_4_9_0_Clk),
    .D(_029_),
    .Q(\memblk.FIFO[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _840_ (.CLK(clknet_4_6_0_Clk),
    .D(_030_),
    .Q(\memblk.FIFO[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _841_ (.CLK(clknet_4_3_0_Clk),
    .D(_031_),
    .Q(\memblk.FIFO[2][31] ));
 sky130_fd_sc_hd__dfrtp_1 _842_ (.CLK(clknet_4_2_0_Clk),
    .D(_032_),
    .RESET_B(net74),
    .Q(\memblk.wr_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _843_ (.CLK(clknet_4_2_0_Clk),
    .D(_033_),
    .RESET_B(net74),
    .Q(\memblk.wr_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _844_ (.CLK(clknet_4_1_0_Clk),
    .D(_034_),
    .Q(\memblk.FIFO[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _845_ (.CLK(clknet_4_2_0_Clk),
    .D(_035_),
    .Q(\memblk.FIFO[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _846_ (.CLK(clknet_4_0_0_Clk),
    .D(_036_),
    .Q(\memblk.FIFO[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _847_ (.CLK(clknet_4_0_0_Clk),
    .D(_037_),
    .Q(\memblk.FIFO[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _848_ (.CLK(clknet_4_6_0_Clk),
    .D(_038_),
    .Q(\memblk.FIFO[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _849_ (.CLK(clknet_4_1_0_Clk),
    .D(_039_),
    .Q(\memblk.FIFO[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _850_ (.CLK(clknet_4_7_0_Clk),
    .D(_040_),
    .Q(\memblk.FIFO[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _851_ (.CLK(clknet_4_5_0_Clk),
    .D(_041_),
    .Q(\memblk.FIFO[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _852_ (.CLK(clknet_4_5_0_Clk),
    .D(_042_),
    .Q(\memblk.FIFO[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _853_ (.CLK(clknet_4_6_0_Clk),
    .D(_043_),
    .Q(\memblk.FIFO[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _854_ (.CLK(clknet_4_6_0_Clk),
    .D(_044_),
    .Q(\memblk.FIFO[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _855_ (.CLK(clknet_4_7_0_Clk),
    .D(_045_),
    .Q(\memblk.FIFO[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _856_ (.CLK(clknet_4_12_0_Clk),
    .D(_046_),
    .Q(\memblk.FIFO[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _857_ (.CLK(clknet_4_13_0_Clk),
    .D(_047_),
    .Q(\memblk.FIFO[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _858_ (.CLK(clknet_4_15_0_Clk),
    .D(_048_),
    .Q(\memblk.FIFO[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _859_ (.CLK(clknet_4_13_0_Clk),
    .D(_049_),
    .Q(\memblk.FIFO[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _860_ (.CLK(clknet_4_13_0_Clk),
    .D(_050_),
    .Q(\memblk.FIFO[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _861_ (.CLK(clknet_4_15_0_Clk),
    .D(_051_),
    .Q(\memblk.FIFO[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _862_ (.CLK(clknet_4_11_0_Clk),
    .D(_052_),
    .Q(\memblk.FIFO[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _863_ (.CLK(clknet_4_14_0_Clk),
    .D(_053_),
    .Q(\memblk.FIFO[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _864_ (.CLK(clknet_4_14_0_Clk),
    .D(_054_),
    .Q(\memblk.FIFO[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _865_ (.CLK(clknet_4_15_0_Clk),
    .D(_055_),
    .Q(\memblk.FIFO[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _866_ (.CLK(clknet_4_12_0_Clk),
    .D(_056_),
    .Q(\memblk.FIFO[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _867_ (.CLK(clknet_4_11_0_Clk),
    .D(_057_),
    .Q(\memblk.FIFO[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _868_ (.CLK(clknet_4_11_0_Clk),
    .D(_058_),
    .Q(\memblk.FIFO[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _869_ (.CLK(clknet_4_8_0_Clk),
    .D(_059_),
    .Q(\memblk.FIFO[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _870_ (.CLK(clknet_4_10_0_Clk),
    .D(_060_),
    .Q(\memblk.FIFO[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _871_ (.CLK(clknet_4_8_0_Clk),
    .D(_061_),
    .Q(\memblk.FIFO[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _872_ (.CLK(clknet_4_10_0_Clk),
    .D(_062_),
    .Q(\memblk.FIFO[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _873_ (.CLK(clknet_4_9_0_Clk),
    .D(_063_),
    .Q(\memblk.FIFO[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _874_ (.CLK(clknet_4_3_0_Clk),
    .D(_064_),
    .Q(\memblk.FIFO[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _875_ (.CLK(clknet_4_9_0_Clk),
    .D(_065_),
    .Q(\memblk.FIFO[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _876_ (.CLK(clknet_4_1_0_Clk),
    .D(_066_),
    .Q(\memblk.FIFO[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _877_ (.CLK(clknet_4_3_0_Clk),
    .D(_067_),
    .Q(\memblk.FIFO[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _878_ (.CLK(clknet_4_0_0_Clk),
    .D(_068_),
    .Q(\memblk.FIFO[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _879_ (.CLK(clknet_4_0_0_Clk),
    .D(_069_),
    .Q(\memblk.FIFO[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _880_ (.CLK(clknet_4_3_0_Clk),
    .D(_070_),
    .Q(\memblk.FIFO[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _881_ (.CLK(clknet_4_1_0_Clk),
    .D(_071_),
    .Q(\memblk.FIFO[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _882_ (.CLK(clknet_4_7_0_Clk),
    .D(_072_),
    .Q(\memblk.FIFO[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _883_ (.CLK(clknet_4_5_0_Clk),
    .D(_073_),
    .Q(\memblk.FIFO[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _884_ (.CLK(clknet_4_4_0_Clk),
    .D(_074_),
    .Q(\memblk.FIFO[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _885_ (.CLK(clknet_4_4_0_Clk),
    .D(_075_),
    .Q(\memblk.FIFO[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _886_ (.CLK(clknet_4_6_0_Clk),
    .D(_076_),
    .Q(\memblk.FIFO[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _887_ (.CLK(clknet_4_7_0_Clk),
    .D(_077_),
    .Q(\memblk.FIFO[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _888_ (.CLK(clknet_4_6_0_Clk),
    .D(_078_),
    .Q(\memblk.FIFO[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _889_ (.CLK(clknet_4_13_0_Clk),
    .D(_079_),
    .Q(\memblk.FIFO[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _890_ (.CLK(clknet_4_13_0_Clk),
    .D(_080_),
    .Q(\memblk.FIFO[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _891_ (.CLK(clknet_4_13_0_Clk),
    .D(_081_),
    .Q(\memblk.FIFO[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _892_ (.CLK(clknet_4_13_0_Clk),
    .D(_082_),
    .Q(\memblk.FIFO[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _893_ (.CLK(clknet_4_12_0_Clk),
    .D(_083_),
    .Q(\memblk.FIFO[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _894_ (.CLK(clknet_4_11_0_Clk),
    .D(_084_),
    .Q(\memblk.FIFO[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _895_ (.CLK(clknet_4_14_0_Clk),
    .D(_085_),
    .Q(\memblk.FIFO[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _896_ (.CLK(clknet_4_14_0_Clk),
    .D(_086_),
    .Q(\memblk.FIFO[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _897_ (.CLK(clknet_4_15_0_Clk),
    .D(_087_),
    .Q(\memblk.FIFO[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _898_ (.CLK(clknet_4_12_0_Clk),
    .D(_088_),
    .Q(\memblk.FIFO[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _899_ (.CLK(clknet_4_11_0_Clk),
    .D(_089_),
    .Q(\memblk.FIFO[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _900_ (.CLK(clknet_4_11_0_Clk),
    .D(_090_),
    .Q(\memblk.FIFO[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _901_ (.CLK(clknet_4_10_0_Clk),
    .D(_091_),
    .Q(\memblk.FIFO[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _902_ (.CLK(clknet_4_10_0_Clk),
    .D(_092_),
    .Q(\memblk.FIFO[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _903_ (.CLK(clknet_4_10_0_Clk),
    .D(_093_),
    .Q(\memblk.FIFO[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _904_ (.CLK(clknet_4_10_0_Clk),
    .D(_094_),
    .Q(\memblk.FIFO[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _905_ (.CLK(clknet_4_9_0_Clk),
    .D(_095_),
    .Q(\memblk.FIFO[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _906_ (.CLK(clknet_4_6_0_Clk),
    .D(_096_),
    .Q(\memblk.FIFO[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _907_ (.CLK(clknet_4_9_0_Clk),
    .D(_097_),
    .Q(\memblk.FIFO[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _908_ (.CLK(clknet_4_1_0_Clk),
    .D(_098_),
    .Q(\memblk.FIFO[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _909_ (.CLK(clknet_4_2_0_Clk),
    .D(_099_),
    .Q(\memblk.FIFO[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _910_ (.CLK(clknet_4_0_0_Clk),
    .D(_100_),
    .Q(\memblk.FIFO[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _911_ (.CLK(clknet_4_0_0_Clk),
    .D(_101_),
    .Q(\memblk.FIFO[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _912_ (.CLK(clknet_4_1_0_Clk),
    .D(_102_),
    .Q(\memblk.FIFO[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _913_ (.CLK(clknet_4_1_0_Clk),
    .D(_103_),
    .Q(\memblk.FIFO[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _914_ (.CLK(clknet_4_5_0_Clk),
    .D(_104_),
    .Q(\memblk.FIFO[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _915_ (.CLK(clknet_4_5_0_Clk),
    .D(_105_),
    .Q(\memblk.FIFO[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _916_ (.CLK(clknet_4_4_0_Clk),
    .D(_106_),
    .Q(\memblk.FIFO[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _917_ (.CLK(clknet_4_4_0_Clk),
    .D(_107_),
    .Q(\memblk.FIFO[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _918_ (.CLK(clknet_4_4_0_Clk),
    .D(_108_),
    .Q(\memblk.FIFO[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _919_ (.CLK(clknet_4_5_0_Clk),
    .D(_109_),
    .Q(\memblk.FIFO[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _920_ (.CLK(clknet_4_6_0_Clk),
    .D(_110_),
    .Q(\memblk.FIFO[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _921_ (.CLK(clknet_4_7_0_Clk),
    .D(_111_),
    .Q(\memblk.FIFO[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _922_ (.CLK(clknet_4_13_0_Clk),
    .D(_112_),
    .Q(\memblk.FIFO[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _923_ (.CLK(clknet_4_7_0_Clk),
    .D(_113_),
    .Q(\memblk.FIFO[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _924_ (.CLK(clknet_4_13_0_Clk),
    .D(_114_),
    .Q(\memblk.FIFO[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _925_ (.CLK(clknet_4_12_0_Clk),
    .D(_115_),
    .Q(\memblk.FIFO[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _926_ (.CLK(clknet_4_9_0_Clk),
    .D(_116_),
    .Q(\memblk.FIFO[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _927_ (.CLK(clknet_4_14_0_Clk),
    .D(_117_),
    .Q(\memblk.FIFO[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _928_ (.CLK(clknet_4_14_0_Clk),
    .D(_118_),
    .Q(\memblk.FIFO[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _929_ (.CLK(clknet_4_15_0_Clk),
    .D(_119_),
    .Q(\memblk.FIFO[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _930_ (.CLK(clknet_4_12_0_Clk),
    .D(_120_),
    .Q(\memblk.FIFO[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _931_ (.CLK(clknet_4_11_0_Clk),
    .D(_121_),
    .Q(\memblk.FIFO[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _932_ (.CLK(clknet_4_9_0_Clk),
    .D(_122_),
    .Q(\memblk.FIFO[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _933_ (.CLK(clknet_4_8_0_Clk),
    .D(_123_),
    .Q(\memblk.FIFO[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _934_ (.CLK(clknet_4_10_0_Clk),
    .D(_124_),
    .Q(\memblk.FIFO[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _935_ (.CLK(clknet_4_8_0_Clk),
    .D(_125_),
    .Q(\memblk.FIFO[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _936_ (.CLK(clknet_4_10_0_Clk),
    .D(_126_),
    .Q(\memblk.FIFO[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _937_ (.CLK(clknet_4_9_0_Clk),
    .D(_127_),
    .Q(\memblk.FIFO[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _938_ (.CLK(clknet_4_3_0_Clk),
    .D(_128_),
    .Q(\memblk.FIFO[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _939_ (.CLK(clknet_4_3_0_Clk),
    .D(_129_),
    .Q(\memblk.FIFO[3][31] ));
 sky130_fd_sc_hd__dfstp_1 _940_ (.CLK(clknet_4_2_0_Clk),
    .D(_130_),
    .SET_B(net75),
    .Q(net71));
 sky130_fd_sc_hd__dfstp_1 _941_ (.CLK(clknet_4_2_0_Clk),
    .D(_131_),
    .SET_B(net74),
    .Q(net72));
 sky130_fd_sc_hd__dfstp_1 _942_ (.CLK(clknet_4_2_0_Clk),
    .D(_132_),
    .SET_B(net75),
    .Q(net73));
 sky130_fd_sc_hd__dfstp_1 _943_ (.CLK(clknet_4_0_0_Clk),
    .D(_133_),
    .SET_B(net75),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _944_ (.CLK(clknet_4_0_0_Clk),
    .D(_134_),
    .RESET_B(net75),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _945_ (.CLK(clknet_4_2_0_Clk),
    .D(_135_),
    .RESET_B(net75),
    .Q(\fcounter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _946_ (.CLK(clknet_4_8_0_Clk),
    .D(_136_),
    .RESET_B(net74),
    .Q(\fcounter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _947_ (.CLK(clknet_4_8_0_Clk),
    .D(_137_),
    .RESET_B(net74),
    .Q(\fcounter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _948_ (.CLK(clknet_4_2_0_Clk),
    .D(_138_),
    .RESET_B(net74),
    .Q(\memblk.rd_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _949_ (.CLK(clknet_4_3_0_Clk),
    .D(_139_),
    .RESET_B(net36),
    .Q(\memblk.rd_addr[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Clk (.A(Clk),
    .X(clknet_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_0_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_10_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_11_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_12_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_13_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_14_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_15_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_1_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_2_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_3_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_4_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_5_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_6_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_7_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_8_0_Clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_Clk (.A(clknet_0_Clk),
    .X(clknet_4_9_0_Clk));
 sky130_fd_sc_hd__clkinv_1 clkload0 (.A(clknet_4_1_0_Clk));
 sky130_fd_sc_hd__clkinv_1 clkload1 (.A(clknet_4_2_0_Clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_4_11_0_Clk));
 sky130_fd_sc_hd__clkinv_2 clkload11 (.A(clknet_4_12_0_Clk));
 sky130_fd_sc_hd__clkbuf_4 clkload12 (.A(clknet_4_13_0_Clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_4_14_0_Clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload14 (.A(clknet_4_15_0_Clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload2 (.A(clknet_4_3_0_Clk));
 sky130_fd_sc_hd__clkinv_1 clkload3 (.A(clknet_4_4_0_Clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_5_0_Clk));
 sky130_fd_sc_hd__clkinv_1 clkload5 (.A(clknet_4_6_0_Clk));
 sky130_fd_sc_hd__clkinv_2 clkload6 (.A(clknet_4_7_0_Clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload7 (.A(clknet_4_8_0_Clk));
 sky130_fd_sc_hd__clkbuf_4 clkload8 (.A(clknet_4_9_0_Clk));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_4_10_0_Clk));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net36),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\memblk.FIFO[3][15] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\memblk.FIFO[3][8] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\memblk.FIFO[1][15] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\memblk.FIFO[0][0] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\memblk.FIFO[1][1] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\memblk.FIFO[0][5] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\memblk.FIFO[2][26] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\memblk.FIFO[0][16] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\memblk.FIFO[1][27] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\memblk.FIFO[1][29] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\memblk.FIFO[2][8] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\memblk.FIFO[3][21] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\memblk.FIFO[3][0] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\memblk.FIFO[2][17] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\memblk.FIFO[2][2] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\memblk.FIFO[2][7] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\memblk.FIFO[2][31] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\memblk.FIFO[0][25] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\memblk.FIFO[2][19] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\memblk.FIFO[2][1] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\memblk.FIFO[0][29] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\memblk.FIFO[0][14] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\memblk.FIFO[0][13] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\memblk.FIFO[0][9] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\memblk.FIFO[1][3] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\memblk.FIFO[1][16] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\memblk.FIFO[1][30] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\memblk.FIFO[2][28] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\memblk.FIFO[0][3] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\memblk.FIFO[1][25] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\memblk.FIFO[0][18] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\memblk.FIFO[1][31] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\memblk.FIFO[0][28] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\memblk.wr_addr[1] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\memblk.FIFO[3][13] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\memblk.FIFO[3][25] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\memblk.FIFO[1][0] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\memblk.FIFO[1][23] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\memblk.FIFO[3][19] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\memblk.FIFO[1][21] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\memblk.FIFO[3][30] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\memblk.FIFO[3][27] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\memblk.FIFO[2][12] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\memblk.FIFO[3][10] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\memblk.FIFO[3][6] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\memblk.FIFO[3][17] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\memblk.FIFO[3][28] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\memblk.FIFO[3][23] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\memblk.FIFO[3][9] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\memblk.FIFO[2][14] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\memblk.FIFO[2][9] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\memblk.FIFO[1][10] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\memblk.FIFO[3][7] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\memblk.FIFO[0][23] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\memblk.FIFO[0][10] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\memblk.FIFO[2][11] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\memblk.FIFO[3][24] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\memblk.FIFO[3][29] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\memblk.FIFO[1][4] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\memblk.FIFO[0][12] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\memblk.FIFO[2][0] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\memblk.FIFO[2][23] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\memblk.FIFO[2][10] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\memblk.FIFO[3][31] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\memblk.FIFO[0][8] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\memblk.FIFO[3][16] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\memblk.FIFO[2][24] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\memblk.FIFO[3][11] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\memblk.FIFO[3][22] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\memblk.FIFO[0][27] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\memblk.FIFO[0][7] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\memblk.FIFO[2][3] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\memblk.FIFO[2][20] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\memblk.FIFO[2][4] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\memblk.FIFO[3][3] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\memblk.FIFO[2][13] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\memblk.FIFO[1][14] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\memblk.FIFO[3][26] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\memblk.FIFO[3][1] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\memblk.FIFO[0][2] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\memblk.FIFO[3][14] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\memblk.FIFO[3][5] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\memblk.FIFO[1][9] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\memblk.FIFO[0][1] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\memblk.FIFO[2][5] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\memblk.FIFO[3][18] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\memblk.FIFO[1][24] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\memblk.FIFO[1][18] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\memblk.FIFO[0][24] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\memblk.FIFO[0][15] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\memblk.FIFO[2][6] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\memblk.FIFO[1][22] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\memblk.FIFO[0][21] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\memblk.FIFO[2][30] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\memblk.FIFO[1][12] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\memblk.FIFO[0][4] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\memblk.FIFO[3][2] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\memblk.FIFO[3][12] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\memblk.FIFO[2][25] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\memblk.FIFO[2][29] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\memblk.FIFO[1][2] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\memblk.FIFO[1][6] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\memblk.FIFO[0][22] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\memblk.FIFO[1][19] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\memblk.FIFO[1][17] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\memblk.FIFO[1][7] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\memblk.FIFO[1][28] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\memblk.FIFO[3][4] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\memblk.FIFO[2][27] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\memblk.FIFO[0][6] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\memblk.FIFO[2][22] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\memblk.FIFO[0][17] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\memblk.FIFO[1][26] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\memblk.FIFO[0][19] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\memblk.FIFO[1][13] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\memblk.FIFO[1][8] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\memblk.FIFO[0][30] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\memblk.FIFO[2][21] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\memblk.FIFO[3][20] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\memblk.FIFO[1][5] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\memblk.FIFO[0][26] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\memblk.FIFO[2][15] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\memblk.FIFO[0][20] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\memblk.FIFO[0][31] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\memblk.FIFO[0][11] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\memblk.FIFO[2][16] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\memblk.FIFO[1][20] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\memblk.FIFO[1][11] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\memblk.FIFO[2][18] ),
    .X(net174));
 sky130_fd_sc_hd__buf_1 input1 (.A(Data_In[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(Data_In[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(Data_In[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(Data_In[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(Data_In[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(Data_In[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(Data_In[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(Data_In[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(Data_In[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(Data_In[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(Data_In[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(Data_In[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(Data_In[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(Data_In[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(Data_In[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(Data_In[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(Data_In[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(Data_In[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(Data_In[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(Data_In[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(Data_In[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(Data_In[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(Data_In[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(Data_In[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(Data_In[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(Data_In[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(FClrN),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(FInN),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(FOutN),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(RstN),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input4 (.A(Data_In[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(Data_In[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(Data_In[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(Data_In[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(Data_In[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(Data_In[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(F_Data[0]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(F_Data[10]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(F_Data[11]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(F_Data[12]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(F_Data[13]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(F_Data[14]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(F_Data[15]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(F_Data[16]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(F_Data[17]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(F_Data[18]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(F_Data[19]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(F_Data[1]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(F_Data[20]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(F_Data[21]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(F_Data[22]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(F_Data[23]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(F_Data[24]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(F_Data[25]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(F_Data[26]));
 sky130_fd_sc_hd__clkbuf_4 output56 (.A(net56),
    .X(F_Data[27]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(F_Data[28]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(F_Data[29]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(F_Data[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(F_Data[30]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(F_Data[31]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(F_Data[3]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(F_Data[4]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(F_Data[5]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(F_Data[6]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(F_Data[7]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(F_Data[8]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(F_Data[9]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(F_EmptyN));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(F_FirstN));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(F_FullN));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(F_LastN));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(F_SLastN));
endmodule

