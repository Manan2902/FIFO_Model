magic
tech sky130A
magscale 1 2
timestamp 1754069373
<< viali >>
rect 10609 24837 10643 24871
rect 4905 24769 4939 24803
rect 6101 24769 6135 24803
rect 7297 24769 7331 24803
rect 8033 24769 8067 24803
rect 8677 24769 8711 24803
rect 9137 24769 9171 24803
rect 10701 24769 10735 24803
rect 11529 24769 11563 24803
rect 12357 24769 12391 24803
rect 13001 24769 13035 24803
rect 13277 24769 13311 24803
rect 13645 24769 13679 24803
rect 14933 24769 14967 24803
rect 15301 24769 15335 24803
rect 15577 24769 15611 24803
rect 15945 24769 15979 24803
rect 16773 24769 16807 24803
rect 18889 24769 18923 24803
rect 20085 24769 20119 24803
rect 20453 24769 20487 24803
rect 20637 24769 20671 24803
rect 5641 24701 5675 24735
rect 6929 24701 6963 24735
rect 10057 24701 10091 24735
rect 10793 24701 10827 24735
rect 12081 24701 12115 24735
rect 14657 24701 14691 24735
rect 18705 24701 18739 24735
rect 19809 24701 19843 24735
rect 4721 24633 4755 24667
rect 6377 24633 6411 24667
rect 8493 24633 8527 24667
rect 13461 24633 13495 24667
rect 4997 24565 5031 24599
rect 6009 24565 6043 24599
rect 7389 24565 7423 24599
rect 8217 24565 8251 24599
rect 9321 24565 9355 24599
rect 9413 24565 9447 24599
rect 10241 24565 10275 24599
rect 12449 24565 12483 24599
rect 13185 24565 13219 24599
rect 13829 24565 13863 24599
rect 14105 24565 14139 24599
rect 16865 24565 16899 24599
rect 18153 24565 18187 24599
rect 19073 24565 19107 24599
rect 19257 24565 19291 24599
rect 20821 24565 20855 24599
rect 5365 24361 5399 24395
rect 11529 24361 11563 24395
rect 12449 24361 12483 24395
rect 16221 24361 16255 24395
rect 19257 24361 19291 24395
rect 5181 24293 5215 24327
rect 17877 24293 17911 24327
rect 9505 24225 9539 24259
rect 13737 24225 13771 24259
rect 16129 24225 16163 24259
rect 16497 24225 16531 24259
rect 18429 24225 18463 24259
rect 18613 24225 18647 24259
rect 3801 24157 3835 24191
rect 5549 24157 5583 24191
rect 5641 24157 5675 24191
rect 7113 24157 7147 24191
rect 8493 24157 8527 24191
rect 8585 24157 8619 24191
rect 9965 24157 9999 24191
rect 11989 24157 12023 24191
rect 12265 24157 12299 24191
rect 12909 24157 12943 24191
rect 13553 24157 13587 24191
rect 14197 24157 14231 24191
rect 14473 24157 14507 24191
rect 16405 24157 16439 24191
rect 20637 24157 20671 24191
rect 4046 24089 4080 24123
rect 5886 24089 5920 24123
rect 10210 24089 10244 24123
rect 11805 24089 11839 24123
rect 15884 24089 15918 24123
rect 16764 24089 16798 24123
rect 18705 24089 18739 24123
rect 20370 24089 20404 24123
rect 7021 24021 7055 24055
rect 7297 24021 7331 24055
rect 8309 24021 8343 24055
rect 8769 24021 8803 24055
rect 8953 24021 8987 24055
rect 9321 24021 9355 24055
rect 9413 24021 9447 24055
rect 11345 24021 11379 24055
rect 12173 24021 12207 24055
rect 12725 24021 12759 24055
rect 13185 24021 13219 24055
rect 13645 24021 13679 24055
rect 14381 24021 14415 24055
rect 14657 24021 14691 24055
rect 14749 24021 14783 24055
rect 19073 24021 19107 24055
rect 3433 23817 3467 23851
rect 5365 23817 5399 23851
rect 5733 23817 5767 23851
rect 6193 23817 6227 23851
rect 9597 23817 9631 23851
rect 9873 23817 9907 23851
rect 11345 23817 11379 23851
rect 13645 23817 13679 23851
rect 16497 23817 16531 23851
rect 16681 23817 16715 23851
rect 17969 23817 18003 23851
rect 21465 23817 21499 23851
rect 7490 23749 7524 23783
rect 8208 23749 8242 23783
rect 10210 23749 10244 23783
rect 12532 23749 12566 23783
rect 13921 23749 13955 23783
rect 20269 23749 20303 23783
rect 3249 23681 3283 23715
rect 3525 23681 3559 23715
rect 3792 23681 3826 23715
rect 5181 23681 5215 23715
rect 5825 23681 5859 23715
rect 9413 23681 9447 23715
rect 9689 23681 9723 23715
rect 9965 23681 9999 23715
rect 12081 23681 12115 23715
rect 14565 23681 14599 23715
rect 14703 23681 14737 23715
rect 14841 23681 14875 23715
rect 15577 23681 15611 23715
rect 15853 23681 15887 23715
rect 16865 23681 16899 23715
rect 17509 23681 17543 23715
rect 20361 23681 20395 23715
rect 20729 23681 20763 23715
rect 21649 23681 21683 23715
rect 5641 23613 5675 23647
rect 7757 23613 7791 23647
rect 7941 23613 7975 23647
rect 12265 23613 12299 23647
rect 15761 23613 15795 23647
rect 17601 23613 17635 23647
rect 17693 23613 17727 23647
rect 18613 23613 18647 23647
rect 18751 23613 18785 23647
rect 18889 23613 18923 23647
rect 19625 23613 19659 23647
rect 19809 23613 19843 23647
rect 20453 23613 20487 23647
rect 21281 23613 21315 23647
rect 6377 23545 6411 23579
rect 15117 23545 15151 23579
rect 19165 23545 19199 23579
rect 4905 23477 4939 23511
rect 9321 23477 9355 23511
rect 11529 23477 11563 23511
rect 17141 23477 17175 23511
rect 19901 23477 19935 23511
rect 3893 23273 3927 23307
rect 5181 23273 5215 23307
rect 8309 23273 8343 23307
rect 10057 23273 10091 23307
rect 13553 23273 13587 23307
rect 16313 23273 16347 23307
rect 17877 23273 17911 23307
rect 20637 23273 20671 23307
rect 7849 23205 7883 23239
rect 8953 23205 8987 23239
rect 11253 23205 11287 23239
rect 4997 23137 5031 23171
rect 5825 23137 5859 23171
rect 5963 23137 5997 23171
rect 6101 23137 6135 23171
rect 6377 23137 6411 23171
rect 6837 23137 6871 23171
rect 7021 23137 7055 23171
rect 7665 23137 7699 23171
rect 9413 23137 9447 23171
rect 9505 23137 9539 23171
rect 10977 23137 11011 23171
rect 11713 23137 11747 23171
rect 11897 23137 11931 23171
rect 15761 23137 15795 23171
rect 15853 23137 15887 23171
rect 18429 23137 18463 23171
rect 18521 23137 18555 23171
rect 4077 23069 4111 23103
rect 8033 23069 8067 23103
rect 8493 23069 8527 23103
rect 10701 23069 10735 23103
rect 10860 23069 10894 23103
rect 12173 23069 12207 23103
rect 12440 23069 12474 23103
rect 14105 23069 14139 23103
rect 16497 23069 16531 23103
rect 18337 23069 18371 23103
rect 18797 23069 18831 23103
rect 19257 23069 19291 23103
rect 14372 23001 14406 23035
rect 15945 23001 15979 23035
rect 16764 23001 16798 23035
rect 19502 23001 19536 23035
rect 4353 22933 4387 22967
rect 4721 22933 4755 22967
rect 4813 22933 4847 22967
rect 7113 22933 7147 22967
rect 9321 22933 9355 22967
rect 15485 22933 15519 22967
rect 17969 22933 18003 22967
rect 18981 22933 19015 22967
rect 4261 22729 4295 22763
rect 5089 22729 5123 22763
rect 6377 22729 6411 22763
rect 6745 22729 6779 22763
rect 6837 22729 6871 22763
rect 9413 22729 9447 22763
rect 10517 22729 10551 22763
rect 10977 22729 11011 22763
rect 13093 22729 13127 22763
rect 14289 22729 14323 22763
rect 14657 22729 14691 22763
rect 16865 22729 16899 22763
rect 17141 22729 17175 22763
rect 17785 22729 17819 22763
rect 19073 22729 19107 22763
rect 4629 22661 4663 22695
rect 8208 22661 8242 22695
rect 10885 22661 10919 22695
rect 13553 22661 13587 22695
rect 15117 22661 15151 22695
rect 4721 22593 4755 22627
rect 5641 22593 5675 22627
rect 6009 22593 6043 22627
rect 10057 22593 10091 22627
rect 13461 22593 13495 22627
rect 14749 22593 14783 22627
rect 15853 22593 15887 22627
rect 17049 22593 17083 22627
rect 17325 22593 17359 22627
rect 18429 22593 18463 22627
rect 18889 22593 18923 22627
rect 4905 22525 4939 22559
rect 6929 22525 6963 22559
rect 7941 22525 7975 22559
rect 11161 22525 11195 22559
rect 13737 22525 13771 22559
rect 14841 22525 14875 22559
rect 15669 22525 15703 22559
rect 16405 22525 16439 22559
rect 9321 22457 9355 22491
rect 5825 22389 5859 22423
rect 5365 22049 5399 22083
rect 6929 22049 6963 22083
rect 9505 22049 9539 22083
rect 4629 21981 4663 22015
rect 6101 21981 6135 22015
rect 6561 21981 6595 22015
rect 7757 21981 7791 22015
rect 9413 21981 9447 22015
rect 10333 21981 10367 22015
rect 10701 21981 10735 22015
rect 12633 21981 12667 22015
rect 12909 21981 12943 22015
rect 14749 21981 14783 22015
rect 15393 21981 15427 22015
rect 16681 21981 16715 22015
rect 19073 21981 19107 22015
rect 20361 21981 20395 22015
rect 5089 21913 5123 21947
rect 7665 21913 7699 21947
rect 9321 21913 9355 21947
rect 9781 21913 9815 21947
rect 3985 21845 4019 21879
rect 4721 21845 4755 21879
rect 5181 21845 5215 21879
rect 5549 21845 5583 21879
rect 7941 21845 7975 21879
rect 8953 21845 8987 21879
rect 10517 21845 10551 21879
rect 12449 21845 12483 21879
rect 12725 21845 12759 21879
rect 14105 21845 14139 21879
rect 14841 21845 14875 21879
rect 16129 21845 16163 21879
rect 18429 21845 18463 21879
rect 19717 21845 19751 21879
rect 6377 21641 6411 21675
rect 11529 21641 11563 21675
rect 13185 21641 13219 21675
rect 13553 21641 13587 21675
rect 14013 21641 14047 21675
rect 14473 21641 14507 21675
rect 15025 21641 15059 21675
rect 18613 21641 18647 21675
rect 5181 21573 5215 21607
rect 11897 21573 11931 21607
rect 3516 21505 3550 21539
rect 5089 21505 5123 21539
rect 6745 21505 6779 21539
rect 6837 21505 6871 21539
rect 7205 21505 7239 21539
rect 8300 21505 8334 21539
rect 9965 21505 9999 21539
rect 10221 21505 10255 21539
rect 11989 21505 12023 21539
rect 12357 21505 12391 21539
rect 13645 21505 13679 21539
rect 14381 21505 14415 21539
rect 16138 21505 16172 21539
rect 16405 21505 16439 21539
rect 16773 21505 16807 21539
rect 17029 21505 17063 21539
rect 18705 21505 18739 21539
rect 19165 21505 19199 21539
rect 19432 21505 19466 21539
rect 23397 21505 23431 21539
rect 3249 21437 3283 21471
rect 5917 21437 5951 21471
rect 6929 21437 6963 21471
rect 7757 21437 7791 21471
rect 8033 21437 8067 21471
rect 12081 21437 12115 21471
rect 12909 21437 12943 21471
rect 13737 21437 13771 21471
rect 14657 21437 14691 21471
rect 18429 21437 18463 21471
rect 20913 21437 20947 21471
rect 18153 21369 18187 21403
rect 4629 21301 4663 21335
rect 9413 21301 9447 21335
rect 11345 21301 11379 21335
rect 19073 21301 19107 21335
rect 20545 21301 20579 21335
rect 21557 21301 21591 21335
rect 23581 21301 23615 21335
rect 3801 21097 3835 21131
rect 8953 21097 8987 21131
rect 16221 21097 16255 21131
rect 16589 21097 16623 21131
rect 20637 21097 20671 21131
rect 13645 21029 13679 21063
rect 18061 21029 18095 21063
rect 4721 20961 4755 20995
rect 5963 20961 5997 20995
rect 6101 20961 6135 20995
rect 6377 20961 6411 20995
rect 7021 20961 7055 20995
rect 10124 20961 10158 20995
rect 10517 20961 10551 20995
rect 10977 20961 11011 20995
rect 14289 20961 14323 20995
rect 14729 20961 14763 20995
rect 15142 20961 15176 20995
rect 15301 20961 15335 20995
rect 18705 20961 18739 20995
rect 19257 20961 19291 20995
rect 21189 20961 21223 20995
rect 21373 20961 21407 20995
rect 3617 20893 3651 20927
rect 3985 20893 4019 20927
rect 4537 20893 4571 20927
rect 4629 20893 4663 20927
rect 5825 20893 5859 20927
rect 6837 20893 6871 20927
rect 8493 20893 8527 20927
rect 8769 20893 8803 20927
rect 9137 20893 9171 20927
rect 9965 20893 9999 20927
rect 10241 20893 10275 20927
rect 11161 20893 11195 20927
rect 11253 20893 11287 20927
rect 12254 20893 12288 20927
rect 12532 20893 12566 20927
rect 13737 20893 13771 20927
rect 14105 20893 14139 20927
rect 15025 20893 15059 20927
rect 15945 20893 15979 20927
rect 16037 20893 16071 20927
rect 16405 20893 16439 20927
rect 16681 20893 16715 20927
rect 18521 20893 18555 20927
rect 8226 20825 8260 20859
rect 11989 20825 12023 20859
rect 16948 20825 16982 20859
rect 19524 20825 19558 20859
rect 21097 20825 21131 20859
rect 3433 20757 3467 20791
rect 4169 20757 4203 20791
rect 5181 20757 5215 20791
rect 7113 20757 7147 20791
rect 8585 20757 8619 20791
rect 9321 20757 9355 20791
rect 13921 20757 13955 20791
rect 18153 20757 18187 20791
rect 18613 20757 18647 20791
rect 20729 20757 20763 20791
rect 4629 20553 4663 20587
rect 6193 20553 6227 20587
rect 7113 20553 7147 20587
rect 9321 20553 9355 20587
rect 9873 20553 9907 20587
rect 11345 20553 11379 20587
rect 13645 20553 13679 20587
rect 15301 20553 15335 20587
rect 15669 20553 15703 20587
rect 20085 20553 20119 20587
rect 20545 20553 20579 20587
rect 8208 20485 8242 20519
rect 10232 20485 10266 20519
rect 12532 20485 12566 20519
rect 17601 20485 17635 20519
rect 3516 20417 3550 20451
rect 5080 20417 5114 20451
rect 6745 20417 6779 20451
rect 7757 20417 7791 20451
rect 7941 20417 7975 20451
rect 9689 20417 9723 20451
rect 9965 20417 9999 20451
rect 12081 20417 12115 20451
rect 13921 20417 13955 20451
rect 14177 20417 14211 20451
rect 15761 20417 15795 20451
rect 16313 20417 16347 20451
rect 16865 20417 16899 20451
rect 18956 20417 18990 20451
rect 19809 20417 19843 20451
rect 19993 20417 20027 20451
rect 20269 20417 20303 20451
rect 20361 20417 20395 20451
rect 23305 20417 23339 20451
rect 23673 20417 23707 20451
rect 3249 20349 3283 20383
rect 4813 20349 4847 20383
rect 6469 20349 6503 20383
rect 6653 20349 6687 20383
rect 7205 20349 7239 20383
rect 12265 20349 12299 20383
rect 15577 20349 15611 20383
rect 18797 20349 18831 20383
rect 19073 20349 19107 20383
rect 19349 20349 19383 20383
rect 16497 20281 16531 20315
rect 11529 20213 11563 20247
rect 16129 20213 16163 20247
rect 18153 20213 18187 20247
rect 23121 20213 23155 20247
rect 23489 20213 23523 20247
rect 7389 20009 7423 20043
rect 8953 20009 8987 20043
rect 10149 20009 10183 20043
rect 11897 20009 11931 20043
rect 14381 20009 14415 20043
rect 16129 20009 16163 20043
rect 17233 20009 17267 20043
rect 19441 20009 19475 20043
rect 9505 19873 9539 19907
rect 10609 19873 10643 19907
rect 10793 19873 10827 19907
rect 14933 19873 14967 19907
rect 15761 19873 15795 19907
rect 17785 19873 17819 19907
rect 18705 19873 18739 19907
rect 7205 19805 7239 19839
rect 9321 19805 9355 19839
rect 10517 19805 10551 19839
rect 11621 19805 11655 19839
rect 12081 19805 12115 19839
rect 14749 19805 14783 19839
rect 15945 19805 15979 19839
rect 17049 19805 17083 19839
rect 17601 19805 17635 19839
rect 19257 19805 19291 19839
rect 22845 19805 22879 19839
rect 22937 19805 22971 19839
rect 23397 19805 23431 19839
rect 23673 19805 23707 19839
rect 9413 19669 9447 19703
rect 14841 19669 14875 19703
rect 15209 19669 15243 19703
rect 17693 19669 17727 19703
rect 18061 19669 18095 19703
rect 22661 19669 22695 19703
rect 23121 19669 23155 19703
rect 23213 19669 23247 19703
rect 23489 19669 23523 19703
rect 7941 19465 7975 19499
rect 9413 19465 9447 19499
rect 11529 19465 11563 19499
rect 13461 19465 13495 19499
rect 15209 19465 15243 19499
rect 16681 19465 16715 19499
rect 1685 19329 1719 19363
rect 3516 19329 3550 19363
rect 6745 19329 6779 19363
rect 6837 19329 6871 19363
rect 8125 19329 8159 19363
rect 10609 19329 10643 19363
rect 11713 19329 11747 19363
rect 13369 19329 13403 19363
rect 13829 19329 13863 19363
rect 15393 19329 15427 19363
rect 16313 19329 16347 19363
rect 16865 19329 16899 19363
rect 17785 19329 17819 19363
rect 20729 19329 20763 19363
rect 21833 19329 21867 19363
rect 23397 19329 23431 19363
rect 3249 19261 3283 19295
rect 5273 19261 5307 19295
rect 6009 19261 6043 19295
rect 6929 19261 6963 19295
rect 7757 19261 7791 19295
rect 9965 19261 9999 19295
rect 11253 19261 11287 19295
rect 13645 19261 13679 19295
rect 14381 19261 14415 19295
rect 18429 19261 18463 19295
rect 19625 19261 19659 19295
rect 22477 19261 22511 19295
rect 23121 19261 23155 19295
rect 4629 19193 4663 19227
rect 1501 19125 1535 19159
rect 4721 19125 4755 19159
rect 5457 19125 5491 19159
rect 6377 19125 6411 19159
rect 7205 19125 7239 19159
rect 10701 19125 10735 19159
rect 13001 19125 13035 19159
rect 16129 19125 16163 19159
rect 20177 19125 20211 19159
rect 20545 19125 20579 19159
rect 22569 19125 22603 19159
rect 23581 19125 23615 19159
rect 3433 18921 3467 18955
rect 5181 18921 5215 18955
rect 7113 18921 7147 18955
rect 22569 18921 22603 18955
rect 1593 18853 1627 18887
rect 13001 18853 13035 18887
rect 19257 18853 19291 18887
rect 21557 18853 21591 18887
rect 4813 18785 4847 18819
rect 5963 18785 5997 18819
rect 6101 18785 6135 18819
rect 6377 18785 6411 18819
rect 6837 18785 6871 18819
rect 8493 18785 8527 18819
rect 10425 18785 10459 18819
rect 13645 18785 13679 18819
rect 15669 18785 15703 18819
rect 19717 18785 19751 18819
rect 19809 18785 19843 18819
rect 20177 18785 20211 18819
rect 22017 18785 22051 18819
rect 22109 18785 22143 18819
rect 1409 18717 1443 18751
rect 3617 18717 3651 18751
rect 3985 18717 4019 18751
rect 4537 18717 4571 18751
rect 5825 18717 5859 18751
rect 7021 18717 7055 18751
rect 9597 18717 9631 18751
rect 11529 18717 11563 18751
rect 12725 18717 12759 18751
rect 13369 18717 13403 18751
rect 14657 18717 14691 18751
rect 15025 18717 15059 18751
rect 15485 18717 15519 18751
rect 16405 18717 16439 18751
rect 18613 18717 18647 18751
rect 18705 18717 18739 18751
rect 19625 18717 19659 18751
rect 20444 18717 20478 18751
rect 23213 18717 23247 18751
rect 23397 18717 23431 18751
rect 4629 18649 4663 18683
rect 8226 18649 8260 18683
rect 10241 18649 10275 18683
rect 10333 18649 10367 18683
rect 10793 18649 10827 18683
rect 16672 18649 16706 18683
rect 3801 18581 3835 18615
rect 4169 18581 4203 18615
rect 8953 18581 8987 18615
rect 9873 18581 9907 18615
rect 12541 18581 12575 18615
rect 13461 18581 13495 18615
rect 14105 18581 14139 18615
rect 14841 18581 14875 18615
rect 16313 18581 16347 18615
rect 17785 18581 17819 18615
rect 17969 18581 18003 18615
rect 18889 18581 18923 18615
rect 22201 18581 22235 18615
rect 22661 18581 22695 18615
rect 23581 18581 23615 18615
rect 4629 18377 4663 18411
rect 4997 18377 5031 18411
rect 6745 18377 6779 18411
rect 8769 18377 8803 18411
rect 9505 18377 9539 18411
rect 10977 18377 11011 18411
rect 11161 18377 11195 18411
rect 13461 18377 13495 18411
rect 15577 18377 15611 18411
rect 16037 18377 16071 18411
rect 19993 18377 20027 18411
rect 21465 18377 21499 18411
rect 3424 18309 3458 18343
rect 5089 18309 5123 18343
rect 6837 18309 6871 18343
rect 7297 18309 7331 18343
rect 8861 18309 8895 18343
rect 9842 18309 9876 18343
rect 12348 18309 12382 18343
rect 15945 18309 15979 18343
rect 5825 18241 5859 18275
rect 8309 18241 8343 18275
rect 9321 18241 9355 18275
rect 9597 18241 9631 18275
rect 11345 18241 11379 18275
rect 11805 18241 11839 18275
rect 14448 18241 14482 18275
rect 14565 18241 14599 18275
rect 16681 18241 16715 18275
rect 18797 18241 18831 18275
rect 19533 18241 19567 18275
rect 19809 18241 19843 18275
rect 20085 18241 20119 18275
rect 20352 18241 20386 18275
rect 22636 18241 22670 18275
rect 3157 18173 3191 18207
rect 5181 18173 5215 18207
rect 6561 18173 6595 18207
rect 7849 18173 7883 18207
rect 8953 18173 8987 18207
rect 12081 18173 12115 18207
rect 13645 18173 13679 18207
rect 14289 18173 14323 18207
rect 15301 18173 15335 18207
rect 15485 18173 15519 18207
rect 16129 18173 16163 18207
rect 17417 18173 17451 18207
rect 18521 18173 18555 18207
rect 18680 18173 18714 18207
rect 19717 18173 19751 18207
rect 22477 18173 22511 18207
rect 22753 18173 22787 18207
rect 23489 18173 23523 18207
rect 23673 18173 23707 18207
rect 4537 18105 4571 18139
rect 8125 18105 8159 18139
rect 14841 18105 14875 18139
rect 19073 18105 19107 18139
rect 23029 18105 23063 18139
rect 5641 18037 5675 18071
rect 7205 18037 7239 18071
rect 8401 18037 8435 18071
rect 11989 18037 12023 18071
rect 17877 18037 17911 18071
rect 21833 18037 21867 18071
rect 6745 17833 6779 17867
rect 7297 17833 7331 17867
rect 9137 17833 9171 17867
rect 13461 17833 13495 17867
rect 15945 17833 15979 17867
rect 17785 17833 17819 17867
rect 19257 17833 19291 17867
rect 23121 17833 23155 17867
rect 8769 17765 8803 17799
rect 10057 17697 10091 17731
rect 10333 17697 10367 17731
rect 10793 17697 10827 17731
rect 11621 17697 11655 17731
rect 12081 17697 12115 17731
rect 18245 17697 18279 17731
rect 18337 17697 18371 17731
rect 21189 17697 21223 17731
rect 21373 17697 21407 17731
rect 5365 17629 5399 17663
rect 7113 17629 7147 17663
rect 7389 17629 7423 17663
rect 9781 17629 9815 17663
rect 9919 17629 9953 17663
rect 10977 17629 11011 17663
rect 12337 17629 12371 17663
rect 13737 17629 13771 17663
rect 14197 17629 14231 17663
rect 14565 17629 14599 17663
rect 16313 17629 16347 17663
rect 18153 17629 18187 17663
rect 18797 17629 18831 17663
rect 20637 17629 20671 17663
rect 21741 17629 21775 17663
rect 23397 17629 23431 17663
rect 5632 17561 5666 17595
rect 7656 17561 7690 17595
rect 11437 17561 11471 17595
rect 14832 17561 14866 17595
rect 16580 17561 16614 17595
rect 20370 17561 20404 17595
rect 21097 17561 21131 17595
rect 21986 17561 22020 17595
rect 11069 17493 11103 17527
rect 11529 17493 11563 17527
rect 13553 17493 13587 17527
rect 14381 17493 14415 17527
rect 17693 17493 17727 17527
rect 18613 17493 18647 17527
rect 20729 17493 20763 17527
rect 23581 17493 23615 17527
rect 7757 17289 7791 17323
rect 8677 17289 8711 17323
rect 11345 17289 11379 17323
rect 11529 17289 11563 17323
rect 14657 17289 14691 17323
rect 16773 17289 16807 17323
rect 17233 17289 17267 17323
rect 17601 17289 17635 17323
rect 19441 17289 19475 17323
rect 20269 17289 20303 17323
rect 22109 17289 22143 17323
rect 23581 17289 23615 17323
rect 13544 17221 13578 17255
rect 18328 17221 18362 17255
rect 21465 17221 21499 17255
rect 22468 17221 22502 17255
rect 5273 17153 5307 17187
rect 5733 17153 5767 17187
rect 5825 17153 5859 17187
rect 6377 17153 6411 17187
rect 7941 17153 7975 17187
rect 8217 17153 8251 17187
rect 8769 17153 8803 17187
rect 9137 17153 9171 17187
rect 9965 17153 9999 17187
rect 10232 17153 10266 17187
rect 12081 17153 12115 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 13277 17153 13311 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 16957 17153 16991 17187
rect 17693 17153 17727 17187
rect 18061 17153 18095 17187
rect 20085 17153 20119 17187
rect 20453 17153 20487 17187
rect 20729 17153 20763 17187
rect 21925 17153 21959 17187
rect 22201 17153 22235 17187
rect 6009 17085 6043 17119
rect 6929 17085 6963 17119
rect 8953 17085 8987 17119
rect 9689 17085 9723 17119
rect 17785 17085 17819 17119
rect 8309 17017 8343 17051
rect 14749 17017 14783 17051
rect 15669 17017 15703 17051
rect 19533 17017 19567 17051
rect 5089 16949 5123 16983
rect 5365 16949 5399 16983
rect 8033 16949 8067 16983
rect 4629 16745 4663 16779
rect 9689 16745 9723 16779
rect 10241 16745 10275 16779
rect 10793 16745 10827 16779
rect 14105 16745 14139 16779
rect 18981 16745 19015 16779
rect 20729 16745 20763 16779
rect 5825 16677 5859 16711
rect 9229 16677 9263 16711
rect 3985 16609 4019 16643
rect 5411 16609 5445 16643
rect 5549 16609 5583 16643
rect 6469 16609 6503 16643
rect 7389 16609 7423 16643
rect 14565 16609 14599 16643
rect 14657 16609 14691 16643
rect 18337 16609 18371 16643
rect 18521 16609 18555 16643
rect 21281 16609 21315 16643
rect 22201 16609 22235 16643
rect 23489 16609 23523 16643
rect 1685 16541 1719 16575
rect 2237 16541 2271 16575
rect 5273 16541 5307 16575
rect 6285 16541 6319 16575
rect 6745 16541 6779 16575
rect 7656 16541 7690 16575
rect 9413 16541 9447 16575
rect 10425 16541 10459 16575
rect 10977 16541 11011 16575
rect 11805 16541 11839 16575
rect 16773 16541 16807 16575
rect 20637 16541 20671 16575
rect 21097 16541 21131 16575
rect 21833 16541 21867 16575
rect 22477 16541 22511 16575
rect 2504 16473 2538 16507
rect 9781 16473 9815 16507
rect 14473 16473 14507 16507
rect 18613 16473 18647 16507
rect 22385 16473 22419 16507
rect 22937 16473 22971 16507
rect 1501 16405 1535 16439
rect 3617 16405 3651 16439
rect 4537 16405 4571 16439
rect 6561 16405 6595 16439
rect 8769 16405 8803 16439
rect 11621 16405 11655 16439
rect 16129 16405 16163 16439
rect 21189 16405 21223 16439
rect 22845 16405 22879 16439
rect 2421 16201 2455 16235
rect 3893 16201 3927 16235
rect 4445 16201 4479 16235
rect 6193 16201 6227 16235
rect 15945 16201 15979 16235
rect 23213 16201 23247 16235
rect 5080 16133 5114 16167
rect 15853 16133 15887 16167
rect 17601 16133 17635 16167
rect 21833 16133 21867 16167
rect 1409 16065 1443 16099
rect 2237 16065 2271 16099
rect 2513 16065 2547 16099
rect 2780 16065 2814 16099
rect 4353 16065 4387 16099
rect 6745 16065 6779 16099
rect 6837 16065 6871 16099
rect 7205 16065 7239 16099
rect 7757 16065 7791 16099
rect 8217 16065 8251 16099
rect 13093 16065 13127 16099
rect 15393 16065 15427 16099
rect 16865 16065 16899 16099
rect 17693 16065 17727 16099
rect 18061 16065 18095 16099
rect 19993 16065 20027 16099
rect 20453 16065 20487 16099
rect 20913 16065 20947 16099
rect 4629 15997 4663 16031
rect 4813 15997 4847 16031
rect 6929 15997 6963 16031
rect 11253 15997 11287 16031
rect 12541 15997 12575 16031
rect 16129 15997 16163 16031
rect 17785 15997 17819 16031
rect 18613 15997 18647 16031
rect 20545 15997 20579 16031
rect 20637 15997 20671 16031
rect 21465 15997 21499 16031
rect 22569 15997 22603 16031
rect 23305 15997 23339 16031
rect 23397 15997 23431 16031
rect 3985 15929 4019 15963
rect 17233 15929 17267 15963
rect 20085 15929 20119 15963
rect 1593 15861 1627 15895
rect 6377 15861 6411 15895
rect 8033 15861 8067 15895
rect 10701 15861 10735 15895
rect 11897 15861 11931 15895
rect 12909 15861 12943 15895
rect 15209 15861 15243 15895
rect 15485 15861 15519 15895
rect 17049 15861 17083 15895
rect 19809 15861 19843 15895
rect 22845 15861 22879 15895
rect 2881 15657 2915 15691
rect 6193 15657 6227 15691
rect 18705 15657 18739 15691
rect 20729 15657 20763 15691
rect 21097 15657 21131 15691
rect 23673 15657 23707 15691
rect 3801 15589 3835 15623
rect 8401 15589 8435 15623
rect 9781 15589 9815 15623
rect 16221 15589 16255 15623
rect 17785 15589 17819 15623
rect 22293 15589 22327 15623
rect 4261 15521 4295 15555
rect 4445 15521 4479 15555
rect 8953 15521 8987 15555
rect 10977 15521 11011 15555
rect 11161 15521 11195 15555
rect 11897 15521 11931 15555
rect 12357 15521 12391 15555
rect 17223 15521 17257 15555
rect 17509 15521 17543 15555
rect 18429 15521 18463 15555
rect 21741 15521 21775 15555
rect 22753 15521 22787 15555
rect 1409 15453 1443 15487
rect 3065 15453 3099 15487
rect 4813 15453 4847 15487
rect 5080 15453 5114 15487
rect 7665 15453 7699 15487
rect 8585 15453 8619 15487
rect 9965 15453 9999 15487
rect 11713 15453 11747 15487
rect 14841 15453 14875 15487
rect 15108 15453 15142 15487
rect 16313 15453 16347 15487
rect 17392 15453 17426 15487
rect 18245 15453 18279 15487
rect 18521 15453 18555 15487
rect 19349 15453 19383 15487
rect 20821 15453 20855 15487
rect 21900 15453 21934 15487
rect 22017 15453 22051 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 10885 15385 10919 15419
rect 11805 15385 11839 15419
rect 12602 15385 12636 15419
rect 19616 15385 19650 15419
rect 1593 15317 1627 15351
rect 4169 15317 4203 15351
rect 8217 15317 8251 15351
rect 9597 15317 9631 15351
rect 10517 15317 10551 15351
rect 11345 15317 11379 15351
rect 13737 15317 13771 15351
rect 16497 15317 16531 15351
rect 16589 15317 16623 15351
rect 21005 15317 21039 15351
rect 3985 15113 4019 15147
rect 5273 15113 5307 15147
rect 7297 15113 7331 15147
rect 7665 15113 7699 15147
rect 7757 15113 7791 15147
rect 11345 15113 11379 15147
rect 11989 15113 12023 15147
rect 14013 15113 14047 15147
rect 16221 15113 16255 15147
rect 18337 15113 18371 15147
rect 18797 15113 18831 15147
rect 23581 15113 23615 15147
rect 14381 15045 14415 15079
rect 17202 15045 17236 15079
rect 1409 14977 1443 15011
rect 4537 14977 4571 15011
rect 5457 14977 5491 15011
rect 7021 14977 7055 15011
rect 9249 14977 9283 15011
rect 9505 14977 9539 15011
rect 9873 14977 9907 15011
rect 9965 14977 9999 15011
rect 10221 14977 10255 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 12725 14977 12759 15011
rect 13001 14977 13035 15011
rect 14841 14977 14875 15011
rect 15108 14977 15142 15011
rect 16681 14977 16715 15011
rect 19616 14977 19650 15011
rect 21189 14977 21223 15011
rect 22946 14977 22980 15011
rect 23213 14977 23247 15011
rect 23397 14977 23431 15011
rect 3617 14909 3651 14943
rect 7849 14909 7883 14943
rect 12863 14909 12897 14943
rect 13277 14909 13311 14943
rect 13737 14909 13771 14943
rect 13921 14909 13955 14943
rect 14473 14909 14507 14943
rect 14657 14909 14691 14943
rect 16957 14909 16991 14943
rect 18889 14909 18923 14943
rect 18981 14909 19015 14943
rect 19349 14909 19383 14943
rect 21281 14909 21315 14943
rect 21465 14909 21499 14943
rect 8125 14841 8159 14875
rect 18429 14841 18463 14875
rect 20729 14841 20763 14875
rect 1593 14773 1627 14807
rect 2973 14773 3007 14807
rect 7205 14773 7239 14807
rect 9689 14773 9723 14807
rect 11529 14773 11563 14807
rect 12081 14773 12115 14807
rect 16865 14773 16899 14807
rect 20821 14773 20855 14807
rect 21833 14773 21867 14807
rect 7297 14569 7331 14603
rect 9781 14569 9815 14603
rect 10333 14569 10367 14603
rect 11989 14569 12023 14603
rect 13921 14569 13955 14603
rect 14841 14569 14875 14603
rect 15577 14569 15611 14603
rect 18705 14569 18739 14603
rect 19257 14569 19291 14603
rect 19993 14569 20027 14603
rect 21005 14569 21039 14603
rect 23305 14569 23339 14603
rect 2421 14501 2455 14535
rect 3801 14501 3835 14535
rect 15025 14501 15059 14535
rect 2973 14433 3007 14467
rect 4445 14433 4479 14467
rect 9137 14433 9171 14467
rect 9229 14433 9263 14467
rect 10609 14433 10643 14467
rect 14197 14433 14231 14467
rect 16037 14433 16071 14467
rect 16129 14433 16163 14467
rect 17049 14433 17083 14467
rect 17325 14433 17359 14467
rect 19809 14433 19843 14467
rect 21649 14433 21683 14467
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 2789 14365 2823 14399
rect 3617 14365 3651 14399
rect 5181 14365 5215 14399
rect 5733 14365 5767 14399
rect 6193 14365 6227 14399
rect 7113 14365 7147 14399
rect 8410 14365 8444 14399
rect 8677 14365 8711 14399
rect 9965 14365 9999 14399
rect 10517 14365 10551 14399
rect 12541 14365 12575 14399
rect 12808 14365 12842 14399
rect 15209 14365 15243 14399
rect 15301 14365 15335 14399
rect 17581 14365 17615 14399
rect 20177 14365 20211 14399
rect 21925 14365 21959 14399
rect 23397 14365 23431 14399
rect 10876 14297 10910 14331
rect 15945 14297 15979 14331
rect 16405 14297 16439 14331
rect 22170 14297 22204 14331
rect 1501 14229 1535 14263
rect 1961 14229 1995 14263
rect 2881 14229 2915 14263
rect 3433 14229 3467 14263
rect 4169 14229 4203 14263
rect 4261 14229 4295 14263
rect 4629 14229 4663 14263
rect 5549 14229 5583 14263
rect 6009 14229 6043 14263
rect 6561 14229 6595 14263
rect 9321 14229 9355 14263
rect 9689 14229 9723 14263
rect 15485 14229 15519 14263
rect 23581 14229 23615 14263
rect 2973 14025 3007 14059
rect 5089 14025 5123 14059
rect 6561 14025 6595 14059
rect 6929 14025 6963 14059
rect 7021 14025 7055 14059
rect 9321 14025 9355 14059
rect 10517 14025 10551 14059
rect 13829 14025 13863 14059
rect 15209 14025 15243 14059
rect 22569 14025 22603 14059
rect 23397 14025 23431 14059
rect 12541 13957 12575 13991
rect 22201 13957 22235 13991
rect 1593 13889 1627 13923
rect 1860 13889 1894 13923
rect 3249 13889 3283 13923
rect 3516 13889 3550 13923
rect 5181 13889 5215 13923
rect 5549 13889 5583 13923
rect 7389 13889 7423 13923
rect 7573 13889 7607 13923
rect 9229 13889 9263 13923
rect 9505 13889 9539 13923
rect 10701 13889 10735 13923
rect 14933 13889 14967 13923
rect 15393 13889 15427 13923
rect 16681 13889 16715 13923
rect 20177 13889 20211 13923
rect 23581 13889 23615 13923
rect 5273 13821 5307 13855
rect 6101 13821 6135 13855
rect 7205 13821 7239 13855
rect 8309 13821 8343 13855
rect 8426 13821 8460 13855
rect 8585 13821 8619 13855
rect 20821 13821 20855 13855
rect 21373 13821 21407 13855
rect 22017 13821 22051 13855
rect 22109 13821 22143 13855
rect 22661 13821 22695 13855
rect 23213 13821 23247 13855
rect 4629 13753 4663 13787
rect 4721 13753 4755 13787
rect 8033 13753 8067 13787
rect 16865 13753 16899 13787
rect 14381 13685 14415 13719
rect 20729 13685 20763 13719
rect 5641 13481 5675 13515
rect 7297 13481 7331 13515
rect 12633 13481 12667 13515
rect 13645 13481 13679 13515
rect 20821 13481 20855 13515
rect 23305 13481 23339 13515
rect 2881 13413 2915 13447
rect 11069 13413 11103 13447
rect 15393 13413 15427 13447
rect 1501 13345 1535 13379
rect 3617 13345 3651 13379
rect 3801 13345 3835 13379
rect 4445 13345 4479 13379
rect 4838 13345 4872 13379
rect 4997 13345 5031 13379
rect 7941 13345 7975 13379
rect 13277 13345 13311 13379
rect 16037 13345 16071 13379
rect 20453 13345 20487 13379
rect 21189 13345 21223 13379
rect 21373 13345 21407 13379
rect 3985 13277 4019 13311
rect 4721 13277 4755 13311
rect 5917 13277 5951 13311
rect 6184 13277 6218 13311
rect 7757 13277 7791 13311
rect 10885 13277 10919 13311
rect 11161 13277 11195 13311
rect 12357 13277 12391 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 15117 13277 15151 13311
rect 16773 13277 16807 13311
rect 17325 13277 17359 13311
rect 17601 13277 17635 13311
rect 19717 13277 19751 13311
rect 21005 13277 21039 13311
rect 21925 13277 21959 13311
rect 23397 13277 23431 13311
rect 1768 13209 1802 13243
rect 2973 13209 3007 13243
rect 13553 13209 13587 13243
rect 15761 13209 15795 13243
rect 16221 13209 16255 13243
rect 21465 13209 21499 13243
rect 22192 13209 22226 13243
rect 7389 13141 7423 13175
rect 7849 13141 7883 13175
rect 11345 13141 11379 13175
rect 11805 13141 11839 13175
rect 14933 13141 14967 13175
rect 15853 13141 15887 13175
rect 17141 13141 17175 13175
rect 17417 13141 17451 13175
rect 19533 13141 19567 13175
rect 19901 13141 19935 13175
rect 20269 13141 20303 13175
rect 20361 13141 20395 13175
rect 21833 13141 21867 13175
rect 23581 13141 23615 13175
rect 1501 12937 1535 12971
rect 1869 12937 1903 12971
rect 2145 12937 2179 12971
rect 2605 12937 2639 12971
rect 5365 12937 5399 12971
rect 7849 12937 7883 12971
rect 9873 12937 9907 12971
rect 11529 12937 11563 12971
rect 13001 12937 13035 12971
rect 15945 12937 15979 12971
rect 16681 12937 16715 12971
rect 18797 12937 18831 12971
rect 20637 12937 20671 12971
rect 21005 12937 21039 12971
rect 2513 12869 2547 12903
rect 3065 12869 3099 12903
rect 12642 12869 12676 12903
rect 1685 12801 1719 12835
rect 2053 12801 2087 12835
rect 3893 12801 3927 12835
rect 3985 12801 4019 12835
rect 4252 12801 4286 12835
rect 6009 12801 6043 12835
rect 6377 12801 6411 12835
rect 6633 12801 6667 12835
rect 8401 12801 8435 12835
rect 8953 12801 8987 12835
rect 9689 12801 9723 12835
rect 10241 12801 10275 12835
rect 10701 12801 10735 12835
rect 13185 12801 13219 12835
rect 14289 12801 14323 12835
rect 14832 12801 14866 12835
rect 17601 12801 17635 12835
rect 18613 12801 18647 12835
rect 18889 12801 18923 12835
rect 19432 12801 19466 12835
rect 21465 12801 21499 12835
rect 22477 12801 22511 12835
rect 22753 12801 22787 12835
rect 23673 12801 23707 12835
rect 2697 12733 2731 12767
rect 10333 12733 10367 12767
rect 10517 12733 10551 12767
rect 11253 12733 11287 12767
rect 12909 12733 12943 12767
rect 14565 12733 14599 12767
rect 17325 12733 17359 12767
rect 17484 12733 17518 12767
rect 17877 12733 17911 12767
rect 18337 12733 18371 12767
rect 18521 12733 18555 12767
rect 19165 12733 19199 12767
rect 21097 12733 21131 12767
rect 21281 12733 21315 12767
rect 22615 12733 22649 12767
rect 23029 12733 23063 12767
rect 23489 12733 23523 12767
rect 6193 12665 6227 12699
rect 7757 12665 7791 12699
rect 8769 12665 8803 12699
rect 20545 12665 20579 12699
rect 21649 12665 21683 12699
rect 9505 12597 9539 12631
rect 14473 12597 14507 12631
rect 19073 12597 19107 12631
rect 21833 12597 21867 12631
rect 3617 12393 3651 12427
rect 10609 12393 10643 12427
rect 14381 12393 14415 12427
rect 16037 12393 16071 12427
rect 18337 12393 18371 12427
rect 20729 12393 20763 12427
rect 21741 12393 21775 12427
rect 23213 12393 23247 12427
rect 1593 12325 1627 12359
rect 10517 12325 10551 12359
rect 11805 12325 11839 12359
rect 15945 12325 15979 12359
rect 20637 12325 20671 12359
rect 23581 12325 23615 12359
rect 11529 12257 11563 12291
rect 12265 12257 12299 12291
rect 14565 12257 14599 12291
rect 16589 12257 16623 12291
rect 18981 12257 19015 12291
rect 19257 12257 19291 12291
rect 21373 12257 21407 12291
rect 21833 12257 21867 12291
rect 1409 12189 1443 12223
rect 3433 12189 3467 12223
rect 3985 12189 4019 12223
rect 8585 12189 8619 12223
rect 9137 12189 9171 12223
rect 9404 12189 9438 12223
rect 11253 12189 11287 12223
rect 11412 12189 11446 12223
rect 12449 12189 12483 12223
rect 13921 12189 13955 12223
rect 14197 12189 14231 12223
rect 14821 12189 14855 12223
rect 16865 12189 16899 12223
rect 17132 12189 17166 12223
rect 19524 12189 19558 12223
rect 21557 12189 21591 12223
rect 22100 12189 22134 12223
rect 23397 12189 23431 12223
rect 13654 12121 13688 12155
rect 16405 12121 16439 12155
rect 8769 12053 8803 12087
rect 12541 12053 12575 12087
rect 16497 12053 16531 12087
rect 18245 12053 18279 12087
rect 18705 12053 18739 12087
rect 18797 12053 18831 12087
rect 1593 11849 1627 11883
rect 10609 11849 10643 11883
rect 11529 11849 11563 11883
rect 11989 11849 12023 11883
rect 12541 11849 12575 11883
rect 16497 11849 16531 11883
rect 16957 11849 16991 11883
rect 18521 11849 18555 11883
rect 19257 11849 19291 11883
rect 20729 11849 20763 11883
rect 21833 11849 21867 11883
rect 17408 11781 17442 11815
rect 1409 11713 1443 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4537 11713 4571 11747
rect 5457 11713 5491 11747
rect 8309 11713 8343 11747
rect 9137 11713 9171 11747
rect 9404 11713 9438 11747
rect 10977 11713 11011 11747
rect 11897 11713 11931 11747
rect 12633 11713 12667 11747
rect 12817 11713 12851 11747
rect 13084 11713 13118 11747
rect 14657 11713 14691 11747
rect 14749 11713 14783 11747
rect 15117 11713 15151 11747
rect 15945 11713 15979 11747
rect 16773 11713 16807 11747
rect 17141 11713 17175 11747
rect 18613 11713 18647 11747
rect 20913 11713 20947 11747
rect 22201 11713 22235 11747
rect 22293 11713 22327 11747
rect 22753 11713 22787 11747
rect 23305 11713 23339 11747
rect 23673 11713 23707 11747
rect 3525 11645 3559 11679
rect 4353 11645 4387 11679
rect 5089 11645 5123 11679
rect 7481 11645 7515 11679
rect 8493 11645 8527 11679
rect 11069 11645 11103 11679
rect 11161 11645 11195 11679
rect 12173 11645 12207 11679
rect 14841 11645 14875 11679
rect 15669 11645 15703 11679
rect 21097 11645 21131 11679
rect 22477 11645 22511 11679
rect 5273 11577 5307 11611
rect 10517 11577 10551 11611
rect 14197 11577 14231 11611
rect 23489 11577 23523 11611
rect 2881 11509 2915 11543
rect 3709 11509 3743 11543
rect 6837 11509 6871 11543
rect 8125 11509 8159 11543
rect 9045 11509 9079 11543
rect 14289 11509 14323 11543
rect 21649 11509 21683 11543
rect 9965 11305 9999 11339
rect 11805 11305 11839 11339
rect 13001 11305 13035 11339
rect 13369 11305 13403 11339
rect 14197 11305 14231 11339
rect 15301 11305 15335 11339
rect 17233 11305 17267 11339
rect 21097 11305 21131 11339
rect 2421 11237 2455 11271
rect 3617 11237 3651 11271
rect 13645 11237 13679 11271
rect 16589 11237 16623 11271
rect 21189 11237 21223 11271
rect 22017 11237 22051 11271
rect 3065 11169 3099 11203
rect 10609 11169 10643 11203
rect 11437 11169 11471 11203
rect 12449 11169 12483 11203
rect 17877 11169 17911 11203
rect 18705 11169 18739 11203
rect 21741 11169 21775 11203
rect 22569 11169 22603 11203
rect 23397 11169 23431 11203
rect 1685 11101 1719 11135
rect 2053 11101 2087 11135
rect 2329 11101 2363 11135
rect 2789 11101 2823 11135
rect 3433 11101 3467 11135
rect 3808 11101 3842 11135
rect 5457 11101 5491 11135
rect 6929 11101 6963 11135
rect 8493 11101 8527 11135
rect 10333 11101 10367 11135
rect 13185 11101 13219 11135
rect 13461 11101 13495 11135
rect 15117 11101 15151 11135
rect 17601 11101 17635 11135
rect 19717 11101 19751 11135
rect 22385 11101 22419 11135
rect 2881 11033 2915 11067
rect 4046 11033 4080 11067
rect 5724 11033 5758 11067
rect 7174 11033 7208 11067
rect 8953 11033 8987 11067
rect 9689 11033 9723 11067
rect 10425 11033 10459 11067
rect 10793 11033 10827 11067
rect 13829 11033 13863 11067
rect 14289 11033 14323 11067
rect 16405 11033 16439 11067
rect 17693 11033 17727 11067
rect 18153 11033 18187 11067
rect 19984 11033 20018 11067
rect 21557 11033 21591 11067
rect 22845 11033 22879 11067
rect 1501 10965 1535 10999
rect 1869 10965 1903 10999
rect 2145 10965 2179 10999
rect 5181 10965 5215 10999
rect 6837 10965 6871 10999
rect 8309 10965 8343 10999
rect 21649 10965 21683 10999
rect 22477 10965 22511 10999
rect 2881 10761 2915 10795
rect 5181 10761 5215 10795
rect 6929 10761 6963 10795
rect 8953 10761 8987 10795
rect 9413 10761 9447 10795
rect 20821 10761 20855 10795
rect 21373 10761 21407 10795
rect 22109 10761 22143 10795
rect 1768 10693 1802 10727
rect 6193 10693 6227 10727
rect 12817 10693 12851 10727
rect 16129 10693 16163 10727
rect 21281 10693 21315 10727
rect 3065 10625 3099 10659
rect 4261 10625 4295 10659
rect 6377 10625 6411 10659
rect 6745 10625 6779 10659
rect 7665 10625 7699 10659
rect 7803 10625 7837 10659
rect 8861 10625 8895 10659
rect 9321 10625 9355 10659
rect 9965 10625 9999 10659
rect 14841 10625 14875 10659
rect 19708 10625 19742 10659
rect 21925 10625 21959 10659
rect 22457 10625 22491 10659
rect 1501 10557 1535 10591
rect 3341 10557 3375 10591
rect 3525 10557 3559 10591
rect 4378 10557 4412 10591
rect 4537 10557 4571 10591
rect 5365 10557 5399 10591
rect 7941 10557 7975 10591
rect 8217 10557 8251 10591
rect 8677 10557 8711 10591
rect 9505 10557 9539 10591
rect 15117 10557 15151 10591
rect 16681 10557 16715 10591
rect 19441 10557 19475 10591
rect 21557 10557 21591 10591
rect 22201 10557 22235 10591
rect 3985 10489 4019 10523
rect 13001 10489 13035 10523
rect 3249 10421 3283 10455
rect 6561 10421 6595 10455
rect 7021 10421 7055 10455
rect 9873 10421 9907 10455
rect 15025 10421 15059 10455
rect 15761 10421 15795 10455
rect 16037 10421 16071 10455
rect 17325 10421 17359 10455
rect 20913 10421 20947 10455
rect 23581 10421 23615 10455
rect 5641 10217 5675 10251
rect 8769 10217 8803 10251
rect 11989 10217 12023 10251
rect 14105 10217 14139 10251
rect 19809 10217 19843 10251
rect 20085 10217 20119 10251
rect 23029 10217 23063 10251
rect 3801 10149 3835 10183
rect 15301 10149 15335 10183
rect 17785 10149 17819 10183
rect 21925 10149 21959 10183
rect 3065 10081 3099 10115
rect 3617 10081 3651 10115
rect 7021 10081 7055 10115
rect 9505 10081 9539 10115
rect 10241 10081 10275 10115
rect 13737 10081 13771 10115
rect 15025 10081 15059 10115
rect 15761 10081 15795 10115
rect 15945 10081 15979 10115
rect 18429 10081 18463 10115
rect 21511 10081 21545 10115
rect 21649 10081 21683 10115
rect 22385 10081 22419 10115
rect 23581 10081 23615 10115
rect 1501 10013 1535 10047
rect 5181 10013 5215 10047
rect 6754 10013 6788 10047
rect 7113 10013 7147 10047
rect 7389 10013 7423 10047
rect 13553 10013 13587 10047
rect 14749 10013 14783 10047
rect 14887 10013 14921 10047
rect 16037 10013 16071 10047
rect 16405 10013 16439 10047
rect 19993 10013 20027 10047
rect 20269 10013 20303 10047
rect 21373 10013 21407 10047
rect 22569 10013 22603 10047
rect 22661 10013 22695 10047
rect 1768 9945 1802 9979
rect 4914 9945 4948 9979
rect 7634 9945 7668 9979
rect 8953 9945 8987 9979
rect 10517 9945 10551 9979
rect 16672 9945 16706 9979
rect 2881 9877 2915 9911
rect 7297 9877 7331 9911
rect 13185 9877 13219 9911
rect 13645 9877 13679 9911
rect 16221 9877 16255 9911
rect 17877 9877 17911 9911
rect 20729 9877 20763 9911
rect 22845 9877 22879 9911
rect 1961 9673 1995 9707
rect 4077 9673 4111 9707
rect 6193 9673 6227 9707
rect 7389 9673 7423 9707
rect 10517 9673 10551 9707
rect 14289 9673 14323 9707
rect 15393 9673 15427 9707
rect 15761 9673 15795 9707
rect 16497 9673 16531 9707
rect 17141 9673 17175 9707
rect 20821 9673 20855 9707
rect 2789 9605 2823 9639
rect 4537 9605 4571 9639
rect 6837 9605 6871 9639
rect 8217 9605 8251 9639
rect 17049 9605 17083 9639
rect 1409 9537 1443 9571
rect 2145 9537 2179 9571
rect 2881 9537 2915 9571
rect 3249 9537 3283 9571
rect 3893 9537 3927 9571
rect 4445 9537 4479 9571
rect 5825 9537 5859 9571
rect 6745 9537 6779 9571
rect 7757 9537 7791 9571
rect 7849 9537 7883 9571
rect 10149 9537 10183 9571
rect 10425 9537 10459 9571
rect 10609 9537 10643 9571
rect 12357 9537 12391 9571
rect 12633 9537 12667 9571
rect 12909 9537 12943 9571
rect 13165 9537 13199 9571
rect 14381 9537 14415 9571
rect 15853 9537 15887 9571
rect 16313 9537 16347 9571
rect 18521 9537 18555 9571
rect 20269 9537 20303 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 21465 9537 21499 9571
rect 22201 9537 22235 9571
rect 22293 9537 22327 9571
rect 22661 9537 22695 9571
rect 23397 9537 23431 9571
rect 3065 9469 3099 9503
rect 4721 9469 4755 9503
rect 5549 9469 5583 9503
rect 5733 9469 5767 9503
rect 6929 9469 6963 9503
rect 7941 9469 7975 9503
rect 9045 9469 9079 9503
rect 15209 9469 15243 9503
rect 15945 9469 15979 9503
rect 17233 9469 17267 9503
rect 18245 9469 18279 9503
rect 18404 9469 18438 9503
rect 19257 9469 19291 9503
rect 19441 9469 19475 9503
rect 20085 9469 20119 9503
rect 22385 9469 22419 9503
rect 23213 9469 23247 9503
rect 2421 9401 2455 9435
rect 12817 9401 12851 9435
rect 18797 9401 18831 9435
rect 21649 9401 21683 9435
rect 23581 9401 23615 9435
rect 1593 9333 1627 9367
rect 6377 9333 6411 9367
rect 10333 9333 10367 9367
rect 12541 9333 12575 9367
rect 16681 9333 16715 9367
rect 17601 9333 17635 9367
rect 19533 9333 19567 9367
rect 21097 9333 21131 9367
rect 21833 9333 21867 9367
rect 5733 9129 5767 9163
rect 6469 9129 6503 9163
rect 9689 9129 9723 9163
rect 9965 9129 9999 9163
rect 12265 9129 12299 9163
rect 15577 9129 15611 9163
rect 18889 9129 18923 9163
rect 20637 9129 20671 9163
rect 22293 9129 22327 9163
rect 22845 9129 22879 9163
rect 1593 9061 1627 9095
rect 9781 9061 9815 9095
rect 23489 9061 23523 9095
rect 3341 8993 3375 9027
rect 5273 8993 5307 9027
rect 6285 8993 6319 9027
rect 9413 8993 9447 9027
rect 10793 8993 10827 9027
rect 12541 8993 12575 9027
rect 14197 8993 14231 9027
rect 16037 8993 16071 9027
rect 1409 8925 1443 8959
rect 2421 8925 2455 8959
rect 4353 8925 4387 8959
rect 6653 8925 6687 8959
rect 9321 8925 9355 8959
rect 10241 8925 10275 8959
rect 10517 8925 10551 8959
rect 12797 8925 12831 8959
rect 15669 8925 15703 8959
rect 17509 8925 17543 8959
rect 19257 8925 19291 8959
rect 20913 8925 20947 8959
rect 21180 8925 21214 8959
rect 22661 8925 22695 8959
rect 23397 8925 23431 8959
rect 23673 8925 23707 8959
rect 3065 8857 3099 8891
rect 3801 8857 3835 8891
rect 14464 8857 14498 8891
rect 16304 8857 16338 8891
rect 17776 8857 17810 8891
rect 19524 8857 19558 8891
rect 2237 8789 2271 8823
rect 2697 8789 2731 8823
rect 3157 8789 3191 8823
rect 4629 8789 4663 8823
rect 4997 8789 5031 8823
rect 5089 8789 5123 8823
rect 8217 8789 8251 8823
rect 13921 8789 13955 8823
rect 15853 8789 15887 8823
rect 17417 8789 17451 8823
rect 23213 8789 23247 8823
rect 3249 8585 3283 8619
rect 3709 8585 3743 8619
rect 6377 8585 6411 8619
rect 9045 8585 9079 8619
rect 9521 8585 9555 8619
rect 9689 8585 9723 8619
rect 13829 8585 13863 8619
rect 15117 8585 15151 8619
rect 16313 8585 16347 8619
rect 16773 8585 16807 8619
rect 17141 8585 17175 8619
rect 17601 8585 17635 8619
rect 18889 8585 18923 8619
rect 19441 8585 19475 8619
rect 2136 8517 2170 8551
rect 9321 8517 9355 8551
rect 14933 8517 14967 8551
rect 18061 8517 18095 8551
rect 19717 8517 19751 8551
rect 1685 8449 1719 8483
rect 3525 8449 3559 8483
rect 4353 8449 4387 8483
rect 4629 8449 4663 8483
rect 5365 8449 5399 8483
rect 5825 8449 5859 8483
rect 8033 8449 8067 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 10149 8449 10183 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 14473 8449 14507 8483
rect 15301 8449 15335 8483
rect 16497 8449 16531 8483
rect 17233 8449 17267 8483
rect 17969 8449 18003 8483
rect 18797 8449 18831 8483
rect 19257 8449 19291 8483
rect 20453 8449 20487 8483
rect 21097 8449 21131 8483
rect 1869 8381 1903 8415
rect 4491 8381 4525 8415
rect 4905 8381 4939 8415
rect 5549 8381 5583 8415
rect 6929 8381 6963 8415
rect 17325 8381 17359 8415
rect 18153 8381 18187 8415
rect 19073 8381 19107 8415
rect 1501 8313 1535 8347
rect 5641 8313 5675 8347
rect 3341 8245 3375 8279
rect 7849 8245 7883 8279
rect 9505 8245 9539 8279
rect 10149 8245 10183 8279
rect 18429 8245 18463 8279
rect 20545 8245 20579 8279
rect 5825 8041 5859 8075
rect 8125 8041 8159 8075
rect 8309 8041 8343 8075
rect 13093 8041 13127 8075
rect 17693 8041 17727 8075
rect 19257 8041 19291 8075
rect 3249 7973 3283 8007
rect 5733 7973 5767 8007
rect 14657 7973 14691 8007
rect 20269 7973 20303 8007
rect 6469 7905 6503 7939
rect 8401 7905 8435 7939
rect 10425 7905 10459 7939
rect 11897 7905 11931 7939
rect 12541 7905 12575 7939
rect 17785 7905 17819 7939
rect 18429 7905 18463 7939
rect 19717 7905 19751 7939
rect 19809 7905 19843 7939
rect 20453 7905 20487 7939
rect 21741 7905 21775 7939
rect 1869 7837 1903 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 4353 7837 4387 7871
rect 7205 7837 7239 7871
rect 7573 7837 7607 7871
rect 7665 7837 7699 7871
rect 7849 7837 7883 7871
rect 7941 7837 7975 7871
rect 8677 7837 8711 7871
rect 10149 7837 10183 7871
rect 12909 7837 12943 7871
rect 13645 7837 13679 7871
rect 14105 7837 14139 7871
rect 14473 7837 14507 7871
rect 17509 7837 17543 7871
rect 19625 7837 19659 7871
rect 20085 7837 20119 7871
rect 2136 7769 2170 7803
rect 4598 7769 4632 7803
rect 6193 7769 6227 7803
rect 12725 7769 12759 7803
rect 20637 7769 20671 7803
rect 21189 7769 21223 7803
rect 3985 7701 4019 7735
rect 4261 7701 4295 7735
rect 6285 7701 6319 7735
rect 6653 7701 6687 7735
rect 7389 7701 7423 7735
rect 11989 7701 12023 7735
rect 13829 7701 13863 7735
rect 14289 7701 14323 7735
rect 20729 7701 20763 7735
rect 21097 7701 21131 7735
rect 3341 7497 3375 7531
rect 5365 7497 5399 7531
rect 8401 7497 8435 7531
rect 12081 7497 12115 7531
rect 12633 7497 12667 7531
rect 13645 7497 13679 7531
rect 20269 7497 20303 7531
rect 4230 7429 4264 7463
rect 15209 7429 15243 7463
rect 19165 7429 19199 7463
rect 21833 7429 21867 7463
rect 2973 7361 3007 7395
rect 8677 7361 8711 7395
rect 8769 7361 8803 7395
rect 8861 7361 8895 7395
rect 9045 7361 9079 7395
rect 9137 7361 9171 7395
rect 9321 7361 9355 7395
rect 11989 7361 12023 7395
rect 12173 7361 12207 7395
rect 12817 7361 12851 7395
rect 13185 7361 13219 7395
rect 13277 7361 13311 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 17509 7361 17543 7395
rect 18429 7361 18463 7395
rect 19073 7361 19107 7395
rect 21382 7361 21416 7395
rect 23397 7361 23431 7395
rect 2789 7293 2823 7327
rect 2881 7293 2915 7327
rect 3985 7293 4019 7327
rect 6469 7293 6503 7327
rect 6837 7293 6871 7327
rect 13369 7293 13403 7327
rect 13921 7293 13955 7327
rect 14473 7293 14507 7327
rect 16313 7293 16347 7327
rect 17233 7293 17267 7327
rect 18061 7293 18095 7327
rect 19257 7293 19291 7327
rect 20085 7293 20119 7327
rect 21649 7293 21683 7327
rect 22385 7293 22419 7327
rect 8263 7157 8297 7191
rect 9137 7157 9171 7191
rect 13093 7157 13127 7191
rect 13277 7157 13311 7191
rect 15761 7157 15795 7191
rect 16681 7157 16715 7191
rect 18245 7157 18279 7191
rect 18705 7157 18739 7191
rect 19533 7157 19567 7191
rect 23581 7157 23615 7191
rect 3801 6953 3835 6987
rect 8033 6953 8067 6987
rect 9505 6953 9539 6987
rect 11805 6953 11839 6987
rect 12265 6953 12299 6987
rect 12909 6953 12943 6987
rect 4353 6817 4387 6851
rect 6469 6817 6503 6851
rect 8677 6817 8711 6851
rect 9045 6817 9079 6851
rect 9229 6817 9263 6851
rect 9597 6817 9631 6851
rect 10149 6817 10183 6851
rect 15209 6817 15243 6851
rect 16037 6817 16071 6851
rect 18889 6817 18923 6851
rect 19809 6817 19843 6851
rect 20453 6817 20487 6851
rect 20729 6817 20763 6851
rect 20867 6817 20901 6851
rect 21005 6817 21039 6851
rect 6101 6749 6135 6783
rect 8953 6749 8987 6783
rect 9505 6749 9539 6783
rect 10057 6749 10091 6783
rect 11345 6749 11379 6783
rect 12356 6749 12390 6783
rect 12449 6749 12483 6783
rect 15761 6749 15795 6783
rect 18061 6749 18095 6783
rect 18705 6749 18739 6783
rect 19993 6749 20027 6783
rect 21741 6749 21775 6783
rect 21997 6749 22031 6783
rect 9229 6681 9263 6715
rect 11989 6681 12023 6715
rect 12725 6681 12759 6715
rect 12941 6681 12975 6715
rect 15025 6681 15059 6715
rect 16304 6681 16338 6715
rect 18797 6681 18831 6715
rect 19349 6681 19383 6715
rect 7895 6613 7929 6647
rect 8401 6613 8435 6647
rect 8493 6613 8527 6647
rect 9873 6613 9907 6647
rect 11529 6613 11563 6647
rect 11621 6613 11655 6647
rect 11789 6613 11823 6647
rect 13093 6613 13127 6647
rect 14657 6613 14691 6647
rect 15117 6613 15151 6647
rect 15945 6613 15979 6647
rect 17417 6613 17451 6647
rect 17509 6613 17543 6647
rect 18337 6613 18371 6647
rect 21649 6613 21683 6647
rect 23121 6613 23155 6647
rect 8217 6409 8251 6443
rect 15577 6409 15611 6443
rect 15945 6409 15979 6443
rect 16681 6409 16715 6443
rect 19625 6409 19659 6443
rect 21373 6409 21407 6443
rect 21649 6409 21683 6443
rect 11805 6341 11839 6375
rect 17794 6341 17828 6375
rect 8309 6273 8343 6307
rect 8677 6273 8711 6307
rect 9505 6273 9539 6307
rect 13553 6273 13587 6307
rect 13829 6273 13863 6307
rect 14105 6273 14139 6307
rect 14361 6273 14395 6307
rect 18512 6273 18546 6307
rect 19973 6273 20007 6307
rect 21189 6273 21223 6307
rect 21465 6273 21499 6307
rect 22753 6273 22787 6307
rect 23673 6273 23707 6307
rect 8401 6205 8435 6239
rect 9873 6205 9907 6239
rect 11529 6205 11563 6239
rect 16037 6205 16071 6239
rect 16129 6205 16163 6239
rect 18061 6205 18095 6239
rect 18245 6205 18279 6239
rect 19717 6205 19751 6239
rect 13737 6137 13771 6171
rect 15485 6137 15519 6171
rect 21097 6137 21131 6171
rect 23489 6137 23523 6171
rect 11299 6069 11333 6103
rect 13277 6069 13311 6103
rect 14013 6069 14047 6103
rect 22201 6069 22235 6103
rect 9781 5865 9815 5899
rect 9965 5865 9999 5899
rect 12265 5865 12299 5899
rect 18521 5865 18555 5899
rect 18981 5865 19015 5899
rect 20821 5865 20855 5899
rect 16865 5797 16899 5831
rect 5089 5729 5123 5763
rect 14105 5729 14139 5763
rect 16451 5729 16485 5763
rect 16589 5729 16623 5763
rect 17325 5729 17359 5763
rect 19901 5729 19935 5763
rect 21281 5729 21315 5763
rect 21465 5729 21499 5763
rect 4721 5661 4755 5695
rect 9137 5661 9171 5695
rect 9321 5661 9355 5695
rect 9413 5661 9447 5695
rect 9505 5661 9539 5695
rect 10149 5661 10183 5695
rect 12081 5661 12115 5695
rect 12842 5661 12876 5695
rect 14361 5661 14395 5695
rect 16313 5661 16347 5695
rect 17509 5661 17543 5695
rect 18705 5661 18739 5695
rect 18797 5661 18831 5695
rect 20729 5661 20763 5695
rect 21189 5661 21223 5695
rect 6515 5593 6549 5627
rect 6653 5593 6687 5627
rect 6837 5593 6871 5627
rect 11529 5593 11563 5627
rect 12449 5593 12483 5627
rect 12633 5593 12667 5627
rect 7021 5525 7055 5559
rect 12771 5525 12805 5559
rect 15485 5525 15519 5559
rect 15669 5525 15703 5559
rect 5825 5321 5859 5355
rect 15301 5321 15335 5355
rect 16221 5321 16255 5355
rect 16681 5321 16715 5355
rect 17141 5321 17175 5355
rect 7297 5253 7331 5287
rect 5733 5185 5767 5219
rect 6101 5185 6135 5219
rect 6653 5185 6687 5219
rect 7021 5185 7055 5219
rect 7113 5185 7147 5219
rect 7481 5185 7515 5219
rect 7665 5185 7699 5219
rect 8033 5185 8067 5219
rect 8125 5185 8159 5219
rect 8953 5185 8987 5219
rect 15853 5185 15887 5219
rect 16405 5185 16439 5219
rect 17049 5185 17083 5219
rect 20085 5185 20119 5219
rect 5825 5117 5859 5151
rect 6377 5117 6411 5151
rect 6561 5117 6595 5151
rect 6745 5117 6779 5151
rect 6837 5117 6871 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 9229 5117 9263 5151
rect 17325 5117 17359 5151
rect 18153 5117 18187 5151
rect 19901 5117 19935 5151
rect 19993 5117 20027 5151
rect 20545 5117 20579 5151
rect 21097 5117 21131 5151
rect 5641 5049 5675 5083
rect 7481 5049 7515 5083
rect 6009 4981 6043 5015
rect 7297 4981 7331 5015
rect 7757 4981 7791 5015
rect 17509 4981 17543 5015
rect 20453 4981 20487 5015
rect 9689 4777 9723 4811
rect 9873 4777 9907 4811
rect 6561 4641 6595 4675
rect 7113 4641 7147 4675
rect 7205 4641 7239 4675
rect 8033 4641 8067 4675
rect 8953 4641 8987 4675
rect 9438 4641 9472 4675
rect 10241 4641 10275 4675
rect 15669 4641 15703 4675
rect 18429 4641 18463 4675
rect 18613 4641 18647 4675
rect 6377 4573 6411 4607
rect 8217 4573 8251 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 10793 4573 10827 4607
rect 10885 4573 10919 4607
rect 12357 4573 12391 4607
rect 17693 4573 17727 4607
rect 19901 4573 19935 4607
rect 21373 4573 21407 4607
rect 7849 4505 7883 4539
rect 9321 4505 9355 4539
rect 9873 4505 9907 4539
rect 15936 4505 15970 4539
rect 17141 4505 17175 4539
rect 18705 4505 18739 4539
rect 19257 4505 19291 4539
rect 21128 4505 21162 4539
rect 5917 4437 5951 4471
rect 6285 4437 6319 4471
rect 7297 4437 7331 4471
rect 7665 4437 7699 4471
rect 9229 4437 9263 4471
rect 9597 4437 9631 4471
rect 10609 4437 10643 4471
rect 12449 4437 12483 4471
rect 17049 4437 17083 4471
rect 19073 4437 19107 4471
rect 19993 4437 20027 4471
rect 6469 4233 6503 4267
rect 7481 4233 7515 4267
rect 10241 4233 10275 4267
rect 10517 4233 10551 4267
rect 17141 4233 17175 4267
rect 19165 4233 19199 4267
rect 21281 4233 21315 4267
rect 8769 4165 8803 4199
rect 11161 4165 11195 4199
rect 5733 4097 5767 4131
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 7665 4097 7699 4131
rect 8033 4097 8067 4131
rect 8401 4097 8435 4131
rect 8493 4097 8527 4131
rect 9229 4097 9263 4131
rect 11345 4097 11379 4131
rect 13277 4097 13311 4131
rect 13461 4097 13495 4131
rect 13728 4097 13762 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 18052 4097 18086 4131
rect 19349 4097 19383 4131
rect 20269 4097 20303 4131
rect 20386 4097 20420 4131
rect 21465 4097 21499 4131
rect 7849 4029 7883 4063
rect 9137 4029 9171 4063
rect 10977 4029 11011 4063
rect 11529 4029 11563 4063
rect 13001 4029 13035 4063
rect 15485 4029 15519 4063
rect 16221 4029 16255 4063
rect 17325 4029 17359 4063
rect 17785 4029 17819 4063
rect 19533 4029 19567 4063
rect 20545 4029 20579 4063
rect 22385 4029 22419 4063
rect 8677 3961 8711 3995
rect 9413 3961 9447 3995
rect 9873 3961 9907 3995
rect 10425 3961 10459 3995
rect 10609 3961 10643 3995
rect 14841 3961 14875 3995
rect 17509 3961 17543 3995
rect 19993 3961 20027 3995
rect 5549 3893 5583 3927
rect 8493 3893 8527 3927
rect 9229 3893 9263 3927
rect 10241 3893 10275 3927
rect 14933 3893 14967 3927
rect 15669 3893 15703 3927
rect 16681 3893 16715 3927
rect 21189 3893 21223 3927
rect 21833 3893 21867 3927
rect 9137 3689 9171 3723
rect 9873 3689 9907 3723
rect 11161 3689 11195 3723
rect 15025 3689 15059 3723
rect 17233 3689 17267 3723
rect 19441 3689 19475 3723
rect 7389 3621 7423 3655
rect 8033 3621 8067 3655
rect 9505 3621 9539 3655
rect 11713 3621 11747 3655
rect 14197 3621 14231 3655
rect 16497 3621 16531 3655
rect 5273 3553 5307 3587
rect 5549 3553 5583 3587
rect 7021 3553 7055 3587
rect 8585 3553 8619 3587
rect 8769 3553 8803 3587
rect 9321 3553 9355 3587
rect 10241 3553 10275 3587
rect 10425 3553 10459 3587
rect 13461 3553 13495 3587
rect 14749 3553 14783 3587
rect 16104 3553 16138 3587
rect 16957 3553 16991 3587
rect 17141 3553 17175 3587
rect 7665 3485 7699 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9413 3485 9447 3519
rect 11529 3485 11563 3519
rect 13921 3485 13955 3519
rect 14565 3485 14599 3519
rect 15209 3485 15243 3519
rect 15945 3485 15979 3519
rect 16221 3485 16255 3519
rect 18613 3485 18647 3519
rect 18889 3485 18923 3519
rect 20821 3485 20855 3519
rect 21465 3485 21499 3519
rect 21833 3485 21867 3519
rect 22109 3485 22143 3519
rect 7205 3417 7239 3451
rect 8033 3417 8067 3451
rect 9873 3417 9907 3451
rect 10517 3417 10551 3451
rect 11161 3417 11195 3451
rect 13185 3417 13219 3451
rect 14657 3417 14691 3451
rect 18346 3417 18380 3451
rect 20576 3417 20610 3451
rect 7481 3349 7515 3383
rect 8493 3349 8527 3383
rect 10057 3349 10091 3383
rect 10885 3349 10919 3383
rect 10977 3349 11011 3383
rect 13737 3349 13771 3383
rect 15301 3349 15335 3383
rect 18705 3349 18739 3383
rect 20913 3349 20947 3383
rect 21649 3349 21683 3383
rect 21925 3349 21959 3383
rect 8401 3145 8435 3179
rect 9597 3145 9631 3179
rect 10425 3145 10459 3179
rect 11713 3145 11747 3179
rect 14841 3145 14875 3179
rect 14933 3145 14967 3179
rect 15393 3145 15427 3179
rect 15945 3145 15979 3179
rect 16957 3145 16991 3179
rect 17049 3145 17083 3179
rect 17417 3145 17451 3179
rect 19717 3145 19751 3179
rect 20453 3145 20487 3179
rect 20821 3145 20855 3179
rect 6929 3077 6963 3111
rect 10701 3077 10735 3111
rect 15301 3077 15335 3111
rect 18052 3077 18086 3111
rect 19625 3077 19659 3111
rect 20361 3077 20395 3111
rect 6653 3009 6687 3043
rect 9781 3009 9815 3043
rect 10885 3009 10919 3043
rect 10977 3009 11011 3043
rect 11529 3009 11563 3043
rect 13461 3009 13495 3043
rect 13728 3009 13762 3043
rect 15761 3009 15795 3043
rect 17693 3009 17727 3043
rect 17785 3009 17819 3043
rect 15577 2941 15611 2975
rect 16865 2941 16899 2975
rect 19809 2941 19843 2975
rect 20177 2941 20211 2975
rect 10057 2873 10091 2907
rect 11161 2873 11195 2907
rect 19165 2873 19199 2907
rect 10425 2805 10459 2839
rect 10609 2805 10643 2839
rect 10701 2805 10735 2839
rect 17509 2805 17543 2839
rect 19257 2805 19291 2839
rect 6101 2601 6135 2635
rect 10793 2601 10827 2635
rect 11069 2601 11103 2635
rect 14473 2601 14507 2635
rect 15761 2601 15795 2635
rect 16405 2601 16439 2635
rect 18153 2601 18187 2635
rect 19625 2601 19659 2635
rect 11897 2533 11931 2567
rect 9413 2465 9447 2499
rect 5917 2397 5951 2431
rect 6653 2397 6687 2431
rect 7573 2397 7607 2431
rect 8125 2397 8159 2431
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 10609 2397 10643 2431
rect 10885 2397 10919 2431
rect 11713 2397 11747 2431
rect 12725 2397 12759 2431
rect 14289 2397 14323 2431
rect 15025 2397 15059 2431
rect 15577 2397 15611 2431
rect 16221 2397 16255 2431
rect 17233 2397 17267 2431
rect 18337 2397 18371 2431
rect 19441 2397 19475 2431
rect 21925 2397 21959 2431
rect 7205 2329 7239 2363
rect 7757 2329 7791 2363
rect 10057 2329 10091 2363
rect 10425 2329 10459 2363
rect 12357 2329 12391 2363
rect 16865 2329 16899 2363
rect 17509 2329 17543 2363
rect 17877 2329 17911 2363
rect 6745 2261 6779 2295
rect 8401 2261 8435 2295
rect 15117 2261 15151 2295
rect 22017 2261 22051 2295
<< metal1 >>
rect 1104 25050 24164 25072
rect 1104 24998 2850 25050
rect 2902 24998 2914 25050
rect 2966 24998 2978 25050
rect 3030 24998 3042 25050
rect 3094 24998 3106 25050
rect 3158 24998 5850 25050
rect 5902 24998 5914 25050
rect 5966 24998 5978 25050
rect 6030 24998 6042 25050
rect 6094 24998 6106 25050
rect 6158 24998 8850 25050
rect 8902 24998 8914 25050
rect 8966 24998 8978 25050
rect 9030 24998 9042 25050
rect 9094 24998 9106 25050
rect 9158 24998 11850 25050
rect 11902 24998 11914 25050
rect 11966 24998 11978 25050
rect 12030 24998 12042 25050
rect 12094 24998 12106 25050
rect 12158 24998 14850 25050
rect 14902 24998 14914 25050
rect 14966 24998 14978 25050
rect 15030 24998 15042 25050
rect 15094 24998 15106 25050
rect 15158 24998 17850 25050
rect 17902 24998 17914 25050
rect 17966 24998 17978 25050
rect 18030 24998 18042 25050
rect 18094 24998 18106 25050
rect 18158 24998 20850 25050
rect 20902 24998 20914 25050
rect 20966 24998 20978 25050
rect 21030 24998 21042 25050
rect 21094 24998 21106 25050
rect 21158 24998 23850 25050
rect 23902 24998 23914 25050
rect 23966 24998 23978 25050
rect 24030 24998 24042 25050
rect 24094 24998 24106 25050
rect 24158 24998 24164 25050
rect 1104 24976 24164 24998
rect 9306 24828 9312 24880
rect 9364 24868 9370 24880
rect 10597 24871 10655 24877
rect 10597 24868 10609 24871
rect 9364 24840 10609 24868
rect 9364 24828 9370 24840
rect 10597 24837 10609 24840
rect 10643 24837 10655 24871
rect 10597 24831 10655 24837
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24800 4951 24803
rect 5166 24800 5172 24812
rect 4939 24772 5172 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5166 24760 5172 24772
rect 5224 24760 5230 24812
rect 6089 24803 6147 24809
rect 6089 24769 6101 24803
rect 6135 24800 6147 24803
rect 6135 24772 7144 24800
rect 6135 24769 6147 24772
rect 6089 24763 6147 24769
rect 5626 24692 5632 24744
rect 5684 24692 5690 24744
rect 6546 24692 6552 24744
rect 6604 24732 6610 24744
rect 6917 24735 6975 24741
rect 6917 24732 6929 24735
rect 6604 24704 6929 24732
rect 6604 24692 6610 24704
rect 6917 24701 6929 24704
rect 6963 24701 6975 24735
rect 7116 24732 7144 24772
rect 7190 24760 7196 24812
rect 7248 24800 7254 24812
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 7248 24772 7297 24800
rect 7248 24760 7254 24772
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 8021 24803 8079 24809
rect 8021 24769 8033 24803
rect 8067 24800 8079 24803
rect 8386 24800 8392 24812
rect 8067 24772 8392 24800
rect 8067 24769 8079 24772
rect 8021 24763 8079 24769
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 8665 24803 8723 24809
rect 8665 24769 8677 24803
rect 8711 24769 8723 24803
rect 8665 24763 8723 24769
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24800 9183 24803
rect 9674 24800 9680 24812
rect 9171 24772 9680 24800
rect 9171 24769 9183 24772
rect 9125 24763 9183 24769
rect 7834 24732 7840 24744
rect 7116 24704 7840 24732
rect 6917 24695 6975 24701
rect 7834 24692 7840 24704
rect 7892 24692 7898 24744
rect 8680 24732 8708 24763
rect 9674 24760 9680 24772
rect 9732 24760 9738 24812
rect 10689 24803 10747 24809
rect 9968 24772 10640 24800
rect 9968 24732 9996 24772
rect 8680 24704 9996 24732
rect 10045 24735 10103 24741
rect 10045 24701 10057 24735
rect 10091 24732 10103 24735
rect 10134 24732 10140 24744
rect 10091 24704 10140 24732
rect 10091 24701 10103 24704
rect 10045 24695 10103 24701
rect 10134 24692 10140 24704
rect 10192 24692 10198 24744
rect 4709 24667 4767 24673
rect 4709 24633 4721 24667
rect 4755 24664 4767 24667
rect 5166 24664 5172 24676
rect 4755 24636 5172 24664
rect 4755 24633 4767 24636
rect 4709 24627 4767 24633
rect 5166 24624 5172 24636
rect 5224 24624 5230 24676
rect 5718 24624 5724 24676
rect 5776 24664 5782 24676
rect 6365 24667 6423 24673
rect 6365 24664 6377 24667
rect 5776 24636 6377 24664
rect 5776 24624 5782 24636
rect 6365 24633 6377 24636
rect 6411 24633 6423 24667
rect 6365 24627 6423 24633
rect 8481 24667 8539 24673
rect 8481 24633 8493 24667
rect 8527 24664 8539 24667
rect 10318 24664 10324 24676
rect 8527 24636 10324 24664
rect 8527 24633 8539 24636
rect 8481 24627 8539 24633
rect 10318 24624 10324 24636
rect 10376 24624 10382 24676
rect 10612 24664 10640 24772
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 10735 24772 11529 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24800 12403 24803
rect 12434 24800 12440 24812
rect 12391 24772 12440 24800
rect 12391 24769 12403 24772
rect 12345 24763 12403 24769
rect 12434 24760 12440 24772
rect 12492 24760 12498 24812
rect 12894 24760 12900 24812
rect 12952 24800 12958 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12952 24772 13001 24800
rect 12952 24760 12958 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24769 13323 24803
rect 13265 24763 13323 24769
rect 10778 24692 10784 24744
rect 10836 24692 10842 24744
rect 11422 24692 11428 24744
rect 11480 24732 11486 24744
rect 12069 24735 12127 24741
rect 12069 24732 12081 24735
rect 11480 24704 12081 24732
rect 11480 24692 11486 24704
rect 12069 24701 12081 24704
rect 12115 24701 12127 24735
rect 12069 24695 12127 24701
rect 12250 24692 12256 24744
rect 12308 24732 12314 24744
rect 13280 24732 13308 24763
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13596 24772 13645 24800
rect 13596 24760 13602 24772
rect 13633 24769 13645 24772
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 14734 24760 14740 24812
rect 14792 24800 14798 24812
rect 14921 24803 14979 24809
rect 14921 24800 14933 24803
rect 14792 24772 14933 24800
rect 14792 24760 14798 24772
rect 14921 24769 14933 24772
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 15528 24772 15577 24800
rect 15528 24760 15534 24772
rect 15565 24769 15577 24772
rect 15611 24769 15623 24803
rect 15565 24763 15623 24769
rect 15933 24803 15991 24809
rect 15933 24769 15945 24803
rect 15979 24800 15991 24803
rect 16206 24800 16212 24812
rect 15979 24772 16212 24800
rect 15979 24769 15991 24772
rect 15933 24763 15991 24769
rect 16206 24760 16212 24772
rect 16264 24760 16270 24812
rect 16761 24803 16819 24809
rect 16761 24769 16773 24803
rect 16807 24769 16819 24803
rect 16761 24763 16819 24769
rect 12308 24704 13308 24732
rect 12308 24692 12314 24704
rect 14642 24692 14648 24744
rect 14700 24692 14706 24744
rect 16022 24692 16028 24744
rect 16080 24732 16086 24744
rect 16776 24732 16804 24763
rect 18782 24760 18788 24812
rect 18840 24800 18846 24812
rect 18877 24803 18935 24809
rect 18877 24800 18889 24803
rect 18840 24772 18889 24800
rect 18840 24760 18846 24772
rect 18877 24769 18889 24772
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19392 24772 19932 24800
rect 19392 24760 19398 24772
rect 16080 24704 16804 24732
rect 18693 24735 18751 24741
rect 16080 24692 16086 24704
rect 18693 24701 18705 24735
rect 18739 24732 18751 24735
rect 19058 24732 19064 24744
rect 18739 24704 19064 24732
rect 18739 24701 18751 24704
rect 18693 24695 18751 24701
rect 19058 24692 19064 24704
rect 19116 24692 19122 24744
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 19797 24735 19855 24741
rect 19797 24732 19809 24735
rect 19300 24704 19809 24732
rect 19300 24692 19306 24704
rect 19797 24701 19809 24704
rect 19843 24701 19855 24735
rect 19904 24732 19932 24772
rect 19978 24760 19984 24812
rect 20036 24800 20042 24812
rect 20073 24803 20131 24809
rect 20073 24800 20085 24803
rect 20036 24772 20085 24800
rect 20036 24760 20042 24772
rect 20073 24769 20085 24772
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 20438 24760 20444 24812
rect 20496 24760 20502 24812
rect 20625 24803 20683 24809
rect 20625 24769 20637 24803
rect 20671 24769 20683 24803
rect 20625 24763 20683 24769
rect 20640 24732 20668 24763
rect 19904 24704 20668 24732
rect 19797 24695 19855 24701
rect 11514 24664 11520 24676
rect 10612 24636 11520 24664
rect 11514 24624 11520 24636
rect 11572 24624 11578 24676
rect 12894 24624 12900 24676
rect 12952 24664 12958 24676
rect 13449 24667 13507 24673
rect 13449 24664 13461 24667
rect 12952 24636 13461 24664
rect 12952 24624 12958 24636
rect 13449 24633 13461 24636
rect 13495 24633 13507 24667
rect 13449 24627 13507 24633
rect 4982 24556 4988 24608
rect 5040 24556 5046 24608
rect 5997 24599 6055 24605
rect 5997 24565 6009 24599
rect 6043 24596 6055 24599
rect 6454 24596 6460 24608
rect 6043 24568 6460 24596
rect 6043 24565 6055 24568
rect 5997 24559 6055 24565
rect 6454 24556 6460 24568
rect 6512 24556 6518 24608
rect 7098 24556 7104 24608
rect 7156 24596 7162 24608
rect 7377 24599 7435 24605
rect 7377 24596 7389 24599
rect 7156 24568 7389 24596
rect 7156 24556 7162 24568
rect 7377 24565 7389 24568
rect 7423 24565 7435 24599
rect 7377 24559 7435 24565
rect 8205 24599 8263 24605
rect 8205 24565 8217 24599
rect 8251 24596 8263 24599
rect 8662 24596 8668 24608
rect 8251 24568 8668 24596
rect 8251 24565 8263 24568
rect 8205 24559 8263 24565
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 9306 24556 9312 24608
rect 9364 24556 9370 24608
rect 9398 24556 9404 24608
rect 9456 24556 9462 24608
rect 9490 24556 9496 24608
rect 9548 24596 9554 24608
rect 10229 24599 10287 24605
rect 10229 24596 10241 24599
rect 9548 24568 10241 24596
rect 9548 24556 9554 24568
rect 10229 24565 10241 24568
rect 10275 24565 10287 24599
rect 10229 24559 10287 24565
rect 11606 24556 11612 24608
rect 11664 24596 11670 24608
rect 12437 24599 12495 24605
rect 12437 24596 12449 24599
rect 11664 24568 12449 24596
rect 11664 24556 11670 24568
rect 12437 24565 12449 24568
rect 12483 24565 12495 24599
rect 12437 24559 12495 24565
rect 13173 24599 13231 24605
rect 13173 24565 13185 24599
rect 13219 24596 13231 24599
rect 13262 24596 13268 24608
rect 13219 24568 13268 24596
rect 13219 24565 13231 24568
rect 13173 24559 13231 24565
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 13814 24556 13820 24608
rect 13872 24556 13878 24608
rect 14090 24556 14096 24608
rect 14148 24556 14154 24608
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 16172 24568 16865 24596
rect 16172 24556 16178 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 16853 24559 16911 24565
rect 18141 24599 18199 24605
rect 18141 24565 18153 24599
rect 18187 24596 18199 24599
rect 18322 24596 18328 24608
rect 18187 24568 18328 24596
rect 18187 24565 18199 24568
rect 18141 24559 18199 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 18966 24556 18972 24608
rect 19024 24596 19030 24608
rect 19061 24599 19119 24605
rect 19061 24596 19073 24599
rect 19024 24568 19073 24596
rect 19024 24556 19030 24568
rect 19061 24565 19073 24568
rect 19107 24565 19119 24599
rect 19061 24559 19119 24565
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 19245 24599 19303 24605
rect 19245 24596 19257 24599
rect 19208 24568 19257 24596
rect 19208 24556 19214 24568
rect 19245 24565 19257 24568
rect 19291 24565 19303 24599
rect 19245 24559 19303 24565
rect 20714 24556 20720 24608
rect 20772 24596 20778 24608
rect 20809 24599 20867 24605
rect 20809 24596 20821 24599
rect 20772 24568 20821 24596
rect 20772 24556 20778 24568
rect 20809 24565 20821 24568
rect 20855 24565 20867 24599
rect 20809 24559 20867 24565
rect 1104 24506 24012 24528
rect 1104 24454 1350 24506
rect 1402 24454 1414 24506
rect 1466 24454 1478 24506
rect 1530 24454 1542 24506
rect 1594 24454 1606 24506
rect 1658 24454 4350 24506
rect 4402 24454 4414 24506
rect 4466 24454 4478 24506
rect 4530 24454 4542 24506
rect 4594 24454 4606 24506
rect 4658 24454 7350 24506
rect 7402 24454 7414 24506
rect 7466 24454 7478 24506
rect 7530 24454 7542 24506
rect 7594 24454 7606 24506
rect 7658 24454 10350 24506
rect 10402 24454 10414 24506
rect 10466 24454 10478 24506
rect 10530 24454 10542 24506
rect 10594 24454 10606 24506
rect 10658 24454 13350 24506
rect 13402 24454 13414 24506
rect 13466 24454 13478 24506
rect 13530 24454 13542 24506
rect 13594 24454 13606 24506
rect 13658 24454 16350 24506
rect 16402 24454 16414 24506
rect 16466 24454 16478 24506
rect 16530 24454 16542 24506
rect 16594 24454 16606 24506
rect 16658 24454 19350 24506
rect 19402 24454 19414 24506
rect 19466 24454 19478 24506
rect 19530 24454 19542 24506
rect 19594 24454 19606 24506
rect 19658 24454 22350 24506
rect 22402 24454 22414 24506
rect 22466 24454 22478 24506
rect 22530 24454 22542 24506
rect 22594 24454 22606 24506
rect 22658 24454 24012 24506
rect 1104 24432 24012 24454
rect 5353 24395 5411 24401
rect 5353 24361 5365 24395
rect 5399 24392 5411 24395
rect 6730 24392 6736 24404
rect 5399 24364 6736 24392
rect 5399 24361 5411 24364
rect 5353 24355 5411 24361
rect 6730 24352 6736 24364
rect 6788 24352 6794 24404
rect 10962 24352 10968 24404
rect 11020 24392 11026 24404
rect 11517 24395 11575 24401
rect 11517 24392 11529 24395
rect 11020 24364 11529 24392
rect 11020 24352 11026 24364
rect 11517 24361 11529 24364
rect 11563 24361 11575 24395
rect 11517 24355 11575 24361
rect 12434 24352 12440 24404
rect 12492 24352 12498 24404
rect 16206 24352 16212 24404
rect 16264 24352 16270 24404
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 5169 24327 5227 24333
rect 5169 24293 5181 24327
rect 5215 24324 5227 24327
rect 5626 24324 5632 24336
rect 5215 24296 5632 24324
rect 5215 24293 5227 24296
rect 5169 24287 5227 24293
rect 5626 24284 5632 24296
rect 5684 24284 5690 24336
rect 17865 24327 17923 24333
rect 17865 24293 17877 24327
rect 17911 24324 17923 24327
rect 19058 24324 19064 24336
rect 17911 24296 19064 24324
rect 17911 24293 17923 24296
rect 17865 24287 17923 24293
rect 19058 24284 19064 24296
rect 19116 24284 19122 24336
rect 9214 24216 9220 24268
rect 9272 24256 9278 24268
rect 9493 24259 9551 24265
rect 9493 24256 9505 24259
rect 9272 24228 9505 24256
rect 9272 24216 9278 24228
rect 9493 24225 9505 24228
rect 9539 24225 9551 24259
rect 9493 24219 9551 24225
rect 13722 24216 13728 24268
rect 13780 24216 13786 24268
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 16206 24256 16212 24268
rect 16163 24228 16212 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 16206 24216 16212 24228
rect 16264 24256 16270 24268
rect 16485 24259 16543 24265
rect 16485 24256 16497 24259
rect 16264 24228 16497 24256
rect 16264 24216 16270 24228
rect 16485 24225 16497 24228
rect 16531 24225 16543 24259
rect 16485 24219 16543 24225
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 18288 24228 18429 24256
rect 18288 24216 18294 24228
rect 18417 24225 18429 24228
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24256 18659 24259
rect 19150 24256 19156 24268
rect 18647 24228 19156 24256
rect 18647 24225 18659 24228
rect 18601 24219 18659 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 3510 24148 3516 24200
rect 3568 24188 3574 24200
rect 3789 24191 3847 24197
rect 3789 24188 3801 24191
rect 3568 24160 3801 24188
rect 3568 24148 3574 24160
rect 3789 24157 3801 24160
rect 3835 24188 3847 24191
rect 3835 24160 5028 24188
rect 3835 24157 3847 24160
rect 3789 24151 3847 24157
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 4034 24123 4092 24129
rect 4034 24120 4046 24123
rect 3476 24092 4046 24120
rect 3476 24080 3482 24092
rect 4034 24089 4046 24092
rect 4080 24089 4092 24123
rect 5000 24120 5028 24160
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24188 5687 24191
rect 5675 24160 6914 24188
rect 5675 24157 5687 24160
rect 5629 24151 5687 24157
rect 5644 24120 5672 24151
rect 5874 24123 5932 24129
rect 5874 24120 5886 24123
rect 5000 24092 5672 24120
rect 5736 24092 5886 24120
rect 4034 24083 4092 24089
rect 5442 24012 5448 24064
rect 5500 24052 5506 24064
rect 5736 24052 5764 24092
rect 5874 24089 5886 24092
rect 5920 24089 5932 24123
rect 6886 24120 6914 24160
rect 7098 24148 7104 24200
rect 7156 24148 7162 24200
rect 8481 24191 8539 24197
rect 8481 24157 8493 24191
rect 8527 24157 8539 24191
rect 8481 24151 8539 24157
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24188 8631 24191
rect 8754 24188 8760 24200
rect 8619 24160 8760 24188
rect 8619 24157 8631 24160
rect 8573 24151 8631 24157
rect 7926 24120 7932 24132
rect 6886 24092 7932 24120
rect 5874 24083 5932 24089
rect 7926 24080 7932 24092
rect 7984 24080 7990 24132
rect 8496 24120 8524 24151
rect 8754 24148 8760 24160
rect 8812 24148 8818 24200
rect 9306 24148 9312 24200
rect 9364 24188 9370 24200
rect 9364 24160 9444 24188
rect 9364 24148 9370 24160
rect 8496 24092 8984 24120
rect 5500 24024 5764 24052
rect 5500 24012 5506 24024
rect 7006 24012 7012 24064
rect 7064 24012 7070 24064
rect 7282 24012 7288 24064
rect 7340 24012 7346 24064
rect 8297 24055 8355 24061
rect 8297 24021 8309 24055
rect 8343 24052 8355 24055
rect 8386 24052 8392 24064
rect 8343 24024 8392 24052
rect 8343 24021 8355 24024
rect 8297 24015 8355 24021
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 8754 24012 8760 24064
rect 8812 24012 8818 24064
rect 8956 24061 8984 24092
rect 8941 24055 8999 24061
rect 8941 24021 8953 24055
rect 8987 24021 8999 24055
rect 8941 24015 8999 24021
rect 9306 24012 9312 24064
rect 9364 24012 9370 24064
rect 9416 24061 9444 24160
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 11977 24191 12035 24197
rect 11977 24157 11989 24191
rect 12023 24157 12035 24191
rect 11977 24151 12035 24157
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 10198 24123 10256 24129
rect 10198 24120 10210 24123
rect 9916 24092 10210 24120
rect 9916 24080 9922 24092
rect 10198 24089 10210 24092
rect 10244 24089 10256 24123
rect 10198 24083 10256 24089
rect 11698 24080 11704 24132
rect 11756 24120 11762 24132
rect 11793 24123 11851 24129
rect 11793 24120 11805 24123
rect 11756 24092 11805 24120
rect 11756 24080 11762 24092
rect 11793 24089 11805 24092
rect 11839 24089 11851 24123
rect 11992 24120 12020 24151
rect 12250 24148 12256 24200
rect 12308 24148 12314 24200
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24188 12955 24191
rect 13541 24191 13599 24197
rect 12943 24160 13216 24188
rect 12943 24157 12955 24160
rect 12897 24151 12955 24157
rect 13078 24120 13084 24132
rect 11992 24092 13084 24120
rect 11793 24083 11851 24089
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 9401 24055 9459 24061
rect 9401 24021 9413 24055
rect 9447 24052 9459 24055
rect 9582 24052 9588 24064
rect 9447 24024 9588 24052
rect 9447 24021 9459 24024
rect 9401 24015 9459 24021
rect 9582 24012 9588 24024
rect 9640 24012 9646 24064
rect 11330 24012 11336 24064
rect 11388 24012 11394 24064
rect 12161 24055 12219 24061
rect 12161 24021 12173 24055
rect 12207 24052 12219 24055
rect 12526 24052 12532 24064
rect 12207 24024 12532 24052
rect 12207 24021 12219 24024
rect 12161 24015 12219 24021
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 12710 24012 12716 24064
rect 12768 24012 12774 24064
rect 13188 24061 13216 24160
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 14090 24188 14096 24200
rect 13587 24160 14096 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14182 24148 14188 24200
rect 14240 24148 14246 24200
rect 14274 24148 14280 24200
rect 14332 24188 14338 24200
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14332 24160 14473 24188
rect 14332 24148 14338 24160
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 14461 24151 14519 24157
rect 14568 24184 16068 24188
rect 16224 24184 16405 24188
rect 14568 24160 16405 24184
rect 13906 24080 13912 24132
rect 13964 24120 13970 24132
rect 14568 24120 14596 24160
rect 16040 24156 16252 24160
rect 16393 24157 16405 24160
rect 16439 24157 16451 24191
rect 20625 24191 20683 24197
rect 20625 24188 20637 24191
rect 16393 24151 16451 24157
rect 20180 24160 20637 24188
rect 20180 24132 20208 24160
rect 20625 24157 20637 24160
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 13964 24092 14596 24120
rect 15872 24123 15930 24129
rect 13964 24080 13970 24092
rect 15872 24089 15884 24123
rect 15918 24120 15930 24123
rect 16574 24120 16580 24132
rect 15918 24092 16580 24120
rect 15918 24089 15930 24092
rect 15872 24083 15930 24089
rect 16574 24080 16580 24092
rect 16632 24080 16638 24132
rect 16752 24123 16810 24129
rect 16752 24089 16764 24123
rect 16798 24120 16810 24123
rect 16850 24120 16856 24132
rect 16798 24092 16856 24120
rect 16798 24089 16810 24092
rect 16752 24083 16810 24089
rect 16850 24080 16856 24092
rect 16908 24080 16914 24132
rect 18414 24080 18420 24132
rect 18472 24120 18478 24132
rect 18693 24123 18751 24129
rect 18693 24120 18705 24123
rect 18472 24092 18705 24120
rect 18472 24080 18478 24092
rect 18693 24089 18705 24092
rect 18739 24120 18751 24123
rect 18966 24120 18972 24132
rect 18739 24092 18972 24120
rect 18739 24089 18751 24092
rect 18693 24083 18751 24089
rect 18966 24080 18972 24092
rect 19024 24120 19030 24132
rect 19610 24120 19616 24132
rect 19024 24092 19616 24120
rect 19024 24080 19030 24092
rect 19610 24080 19616 24092
rect 19668 24080 19674 24132
rect 20162 24080 20168 24132
rect 20220 24080 20226 24132
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 20358 24123 20416 24129
rect 20358 24120 20370 24123
rect 20312 24092 20370 24120
rect 20312 24080 20318 24092
rect 20358 24089 20370 24092
rect 20404 24089 20416 24123
rect 20358 24083 20416 24089
rect 13173 24055 13231 24061
rect 13173 24021 13185 24055
rect 13219 24021 13231 24055
rect 13173 24015 13231 24021
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 13814 24052 13820 24064
rect 13679 24024 13820 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 14366 24012 14372 24064
rect 14424 24012 14430 24064
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 14608 24024 14657 24052
rect 14608 24012 14614 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 14737 24055 14795 24061
rect 14737 24021 14749 24055
rect 14783 24052 14795 24055
rect 15562 24052 15568 24064
rect 14783 24024 15568 24052
rect 14783 24021 14795 24024
rect 14737 24015 14795 24021
rect 15562 24012 15568 24024
rect 15620 24012 15626 24064
rect 18874 24012 18880 24064
rect 18932 24052 18938 24064
rect 19061 24055 19119 24061
rect 19061 24052 19073 24055
rect 18932 24024 19073 24052
rect 18932 24012 18938 24024
rect 19061 24021 19073 24024
rect 19107 24021 19119 24055
rect 19061 24015 19119 24021
rect 1104 23962 24164 23984
rect 1104 23910 2850 23962
rect 2902 23910 2914 23962
rect 2966 23910 2978 23962
rect 3030 23910 3042 23962
rect 3094 23910 3106 23962
rect 3158 23910 5850 23962
rect 5902 23910 5914 23962
rect 5966 23910 5978 23962
rect 6030 23910 6042 23962
rect 6094 23910 6106 23962
rect 6158 23910 8850 23962
rect 8902 23910 8914 23962
rect 8966 23910 8978 23962
rect 9030 23910 9042 23962
rect 9094 23910 9106 23962
rect 9158 23910 11850 23962
rect 11902 23910 11914 23962
rect 11966 23910 11978 23962
rect 12030 23910 12042 23962
rect 12094 23910 12106 23962
rect 12158 23910 14850 23962
rect 14902 23910 14914 23962
rect 14966 23910 14978 23962
rect 15030 23910 15042 23962
rect 15094 23910 15106 23962
rect 15158 23910 17850 23962
rect 17902 23910 17914 23962
rect 17966 23910 17978 23962
rect 18030 23910 18042 23962
rect 18094 23910 18106 23962
rect 18158 23910 20850 23962
rect 20902 23910 20914 23962
rect 20966 23910 20978 23962
rect 21030 23910 21042 23962
rect 21094 23910 21106 23962
rect 21158 23910 23850 23962
rect 23902 23910 23914 23962
rect 23966 23910 23978 23962
rect 24030 23910 24042 23962
rect 24094 23910 24106 23962
rect 24158 23910 24164 23962
rect 1104 23888 24164 23910
rect 3418 23808 3424 23860
rect 3476 23808 3482 23860
rect 5353 23851 5411 23857
rect 5353 23817 5365 23851
rect 5399 23848 5411 23851
rect 5442 23848 5448 23860
rect 5399 23820 5448 23848
rect 5399 23817 5411 23820
rect 5353 23811 5411 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 5718 23808 5724 23860
rect 5776 23808 5782 23860
rect 6181 23851 6239 23857
rect 6181 23817 6193 23851
rect 6227 23848 6239 23851
rect 7098 23848 7104 23860
rect 6227 23820 7104 23848
rect 6227 23817 6239 23820
rect 6181 23811 6239 23817
rect 7098 23808 7104 23820
rect 7156 23808 7162 23860
rect 9585 23851 9643 23857
rect 9585 23817 9597 23851
rect 9631 23817 9643 23851
rect 9585 23811 9643 23817
rect 4246 23780 4252 23792
rect 3252 23752 4252 23780
rect 3252 23721 3280 23752
rect 4246 23740 4252 23752
rect 4304 23740 4310 23792
rect 7282 23740 7288 23792
rect 7340 23780 7346 23792
rect 7478 23783 7536 23789
rect 7478 23780 7490 23783
rect 7340 23752 7490 23780
rect 7340 23740 7346 23752
rect 7478 23749 7490 23752
rect 7524 23749 7536 23783
rect 7478 23743 7536 23749
rect 8196 23783 8254 23789
rect 8196 23749 8208 23783
rect 8242 23780 8254 23783
rect 8294 23780 8300 23792
rect 8242 23752 8300 23780
rect 8242 23749 8254 23752
rect 8196 23743 8254 23749
rect 8294 23740 8300 23752
rect 8352 23740 8358 23792
rect 9600 23780 9628 23811
rect 9858 23808 9864 23860
rect 9916 23808 9922 23860
rect 11333 23851 11391 23857
rect 11333 23817 11345 23851
rect 11379 23848 11391 23851
rect 11422 23848 11428 23860
rect 11379 23820 11428 23848
rect 11379 23817 11391 23820
rect 11333 23811 11391 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 13633 23851 13691 23857
rect 13633 23817 13645 23851
rect 13679 23848 13691 23851
rect 14642 23848 14648 23860
rect 13679 23820 14648 23848
rect 13679 23817 13691 23820
rect 13633 23811 13691 23817
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 15838 23808 15844 23860
rect 15896 23848 15902 23860
rect 16485 23851 16543 23857
rect 16485 23848 16497 23851
rect 15896 23820 16497 23848
rect 15896 23808 15902 23820
rect 16485 23817 16497 23820
rect 16531 23817 16543 23851
rect 16485 23811 16543 23817
rect 16574 23808 16580 23860
rect 16632 23848 16638 23860
rect 16669 23851 16727 23857
rect 16669 23848 16681 23851
rect 16632 23820 16681 23848
rect 16632 23808 16638 23820
rect 16669 23817 16681 23820
rect 16715 23817 16727 23851
rect 16669 23811 16727 23817
rect 17957 23851 18015 23857
rect 17957 23817 17969 23851
rect 18003 23848 18015 23851
rect 18003 23820 20392 23848
rect 18003 23817 18015 23820
rect 17957 23811 18015 23817
rect 10198 23783 10256 23789
rect 10198 23780 10210 23783
rect 9600 23752 10210 23780
rect 10198 23749 10210 23752
rect 10244 23749 10256 23783
rect 10198 23743 10256 23749
rect 12520 23783 12578 23789
rect 12520 23749 12532 23783
rect 12566 23780 12578 23783
rect 12710 23780 12716 23792
rect 12566 23752 12716 23780
rect 12566 23749 12578 23752
rect 12520 23743 12578 23749
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 13906 23740 13912 23792
rect 13964 23740 13970 23792
rect 19610 23740 19616 23792
rect 19668 23780 19674 23792
rect 20257 23783 20315 23789
rect 20257 23780 20269 23783
rect 19668 23752 20269 23780
rect 19668 23740 19674 23752
rect 20257 23749 20269 23752
rect 20303 23749 20315 23783
rect 20364 23780 20392 23820
rect 20438 23808 20444 23860
rect 20496 23848 20502 23860
rect 21453 23851 21511 23857
rect 21453 23848 21465 23851
rect 20496 23820 21465 23848
rect 20496 23808 20502 23820
rect 21453 23817 21465 23820
rect 21499 23817 21511 23851
rect 21453 23811 21511 23817
rect 20364 23752 21680 23780
rect 20257 23743 20315 23749
rect 3237 23715 3295 23721
rect 3237 23681 3249 23715
rect 3283 23681 3295 23715
rect 3237 23675 3295 23681
rect 3510 23672 3516 23724
rect 3568 23672 3574 23724
rect 3786 23721 3792 23724
rect 3780 23675 3792 23721
rect 3786 23672 3792 23675
rect 3844 23672 3850 23724
rect 5169 23715 5227 23721
rect 5169 23681 5181 23715
rect 5215 23712 5227 23715
rect 5813 23715 5871 23721
rect 5215 23684 5764 23712
rect 5215 23681 5227 23684
rect 5169 23675 5227 23681
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23613 5687 23647
rect 5736 23644 5764 23684
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 6730 23712 6736 23724
rect 5859 23684 6736 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23712 9459 23715
rect 9490 23712 9496 23724
rect 9447 23684 9496 23712
rect 9447 23681 9459 23684
rect 9401 23675 9459 23681
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 9674 23672 9680 23724
rect 9732 23672 9738 23724
rect 9950 23672 9956 23724
rect 10008 23672 10014 23724
rect 10778 23712 10784 23724
rect 10060 23684 10784 23712
rect 6270 23644 6276 23656
rect 5736 23616 6276 23644
rect 5629 23607 5687 23613
rect 5644 23576 5672 23607
rect 6270 23604 6276 23616
rect 6328 23604 6334 23656
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23644 7803 23647
rect 7926 23644 7932 23656
rect 7791 23616 7932 23644
rect 7791 23613 7803 23616
rect 7745 23607 7803 23613
rect 7926 23604 7932 23616
rect 7984 23604 7990 23656
rect 10060 23644 10088 23684
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 11330 23672 11336 23724
rect 11388 23712 11394 23724
rect 11882 23712 11888 23724
rect 11388 23684 11888 23712
rect 11388 23672 11394 23684
rect 11882 23672 11888 23684
rect 11940 23712 11946 23724
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 11940 23684 12081 23712
rect 11940 23672 11946 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 9232 23616 10088 23644
rect 6365 23579 6423 23585
rect 5644 23548 6316 23576
rect 4893 23511 4951 23517
rect 4893 23477 4905 23511
rect 4939 23508 4951 23511
rect 5626 23508 5632 23520
rect 4939 23480 5632 23508
rect 4939 23477 4951 23480
rect 4893 23471 4951 23477
rect 5626 23468 5632 23480
rect 5684 23508 5690 23520
rect 6086 23508 6092 23520
rect 5684 23480 6092 23508
rect 5684 23468 5690 23480
rect 6086 23468 6092 23480
rect 6144 23468 6150 23520
rect 6288 23508 6316 23548
rect 6365 23545 6377 23579
rect 6411 23576 6423 23579
rect 6546 23576 6552 23588
rect 6411 23548 6552 23576
rect 6411 23545 6423 23548
rect 6365 23539 6423 23545
rect 6546 23536 6552 23548
rect 6604 23536 6610 23588
rect 6454 23508 6460 23520
rect 6288 23480 6460 23508
rect 6454 23468 6460 23480
rect 6512 23508 6518 23520
rect 9232 23508 9260 23616
rect 12250 23604 12256 23656
rect 12308 23604 12314 23656
rect 14568 23644 14596 23675
rect 14642 23672 14648 23724
rect 14700 23721 14706 23724
rect 14700 23715 14749 23721
rect 14700 23681 14703 23715
rect 14737 23681 14749 23715
rect 14700 23675 14749 23681
rect 14700 23672 14706 23675
rect 14826 23672 14832 23724
rect 14884 23672 14890 23724
rect 15562 23672 15568 23724
rect 15620 23712 15626 23724
rect 15841 23715 15899 23721
rect 15841 23712 15853 23715
rect 15620 23684 15853 23712
rect 15620 23672 15626 23684
rect 15841 23681 15853 23684
rect 15887 23681 15899 23715
rect 15841 23675 15899 23681
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 21652 23721 21680 23752
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16816 23684 16865 23712
rect 16816 23672 16822 23684
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23712 17555 23715
rect 20349 23715 20407 23721
rect 17543 23684 18092 23712
rect 17543 23681 17555 23684
rect 17497 23675 17555 23681
rect 14200 23616 14596 23644
rect 6512 23480 9260 23508
rect 9309 23511 9367 23517
rect 6512 23468 6518 23480
rect 9309 23477 9321 23511
rect 9355 23508 9367 23511
rect 10134 23508 10140 23520
rect 9355 23480 10140 23508
rect 9355 23477 9367 23480
rect 9309 23471 9367 23477
rect 10134 23468 10140 23480
rect 10192 23508 10198 23520
rect 10870 23508 10876 23520
rect 10192 23480 10876 23508
rect 10192 23468 10198 23480
rect 10870 23468 10876 23480
rect 10928 23468 10934 23520
rect 11514 23468 11520 23520
rect 11572 23468 11578 23520
rect 14200 23508 14228 23616
rect 15746 23604 15752 23656
rect 15804 23604 15810 23656
rect 17586 23604 17592 23656
rect 17644 23604 17650 23656
rect 17678 23604 17684 23656
rect 17736 23604 17742 23656
rect 18064 23644 18092 23684
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 20717 23715 20775 23721
rect 20717 23712 20729 23715
rect 20395 23684 20729 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 20717 23681 20729 23684
rect 20763 23681 20775 23715
rect 20717 23675 20775 23681
rect 21637 23715 21695 23721
rect 21637 23681 21649 23715
rect 21683 23681 21695 23715
rect 21637 23675 21695 23681
rect 18414 23644 18420 23656
rect 18064 23616 18420 23644
rect 18414 23604 18420 23616
rect 18472 23604 18478 23656
rect 18598 23604 18604 23656
rect 18656 23604 18662 23656
rect 18690 23604 18696 23656
rect 18748 23653 18754 23656
rect 18748 23647 18797 23653
rect 18748 23613 18751 23647
rect 18785 23613 18797 23647
rect 18748 23607 18797 23613
rect 18877 23647 18935 23653
rect 18877 23613 18889 23647
rect 18923 23644 18935 23647
rect 19058 23644 19064 23656
rect 18923 23616 19064 23644
rect 18923 23613 18935 23616
rect 18877 23607 18935 23613
rect 18748 23604 18754 23607
rect 19058 23604 19064 23616
rect 19116 23604 19122 23656
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 19300 23616 19625 23644
rect 19300 23604 19306 23616
rect 19613 23613 19625 23616
rect 19659 23613 19671 23647
rect 19613 23607 19671 23613
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23644 19855 23647
rect 19978 23644 19984 23656
rect 19843 23616 19984 23644
rect 19843 23613 19855 23616
rect 19797 23607 19855 23613
rect 19978 23604 19984 23616
rect 20036 23604 20042 23656
rect 20438 23604 20444 23656
rect 20496 23604 20502 23656
rect 21269 23647 21327 23653
rect 21269 23613 21281 23647
rect 21315 23613 21327 23647
rect 21269 23607 21327 23613
rect 15102 23536 15108 23588
rect 15160 23536 15166 23588
rect 15488 23548 18276 23576
rect 15488 23520 15516 23548
rect 15470 23508 15476 23520
rect 14200 23480 15476 23508
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 17129 23511 17187 23517
rect 17129 23477 17141 23511
rect 17175 23508 17187 23511
rect 17310 23508 17316 23520
rect 17175 23480 17316 23508
rect 17175 23477 17187 23480
rect 17129 23471 17187 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 18248 23508 18276 23548
rect 19150 23536 19156 23588
rect 19208 23536 19214 23588
rect 19996 23576 20024 23604
rect 21284 23576 21312 23607
rect 19996 23548 21312 23576
rect 18598 23508 18604 23520
rect 18248 23480 18604 23508
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 19886 23468 19892 23520
rect 19944 23468 19950 23520
rect 1104 23418 24012 23440
rect 1104 23366 1350 23418
rect 1402 23366 1414 23418
rect 1466 23366 1478 23418
rect 1530 23366 1542 23418
rect 1594 23366 1606 23418
rect 1658 23366 4350 23418
rect 4402 23366 4414 23418
rect 4466 23366 4478 23418
rect 4530 23366 4542 23418
rect 4594 23366 4606 23418
rect 4658 23366 7350 23418
rect 7402 23366 7414 23418
rect 7466 23366 7478 23418
rect 7530 23366 7542 23418
rect 7594 23366 7606 23418
rect 7658 23366 10350 23418
rect 10402 23366 10414 23418
rect 10466 23366 10478 23418
rect 10530 23366 10542 23418
rect 10594 23366 10606 23418
rect 10658 23366 13350 23418
rect 13402 23366 13414 23418
rect 13466 23366 13478 23418
rect 13530 23366 13542 23418
rect 13594 23366 13606 23418
rect 13658 23366 16350 23418
rect 16402 23366 16414 23418
rect 16466 23366 16478 23418
rect 16530 23366 16542 23418
rect 16594 23366 16606 23418
rect 16658 23366 19350 23418
rect 19402 23366 19414 23418
rect 19466 23366 19478 23418
rect 19530 23366 19542 23418
rect 19594 23366 19606 23418
rect 19658 23366 22350 23418
rect 22402 23366 22414 23418
rect 22466 23366 22478 23418
rect 22530 23366 22542 23418
rect 22594 23366 22606 23418
rect 22658 23366 24012 23418
rect 1104 23344 24012 23366
rect 3786 23264 3792 23316
rect 3844 23304 3850 23316
rect 3881 23307 3939 23313
rect 3881 23304 3893 23307
rect 3844 23276 3893 23304
rect 3844 23264 3850 23276
rect 3881 23273 3893 23276
rect 3927 23273 3939 23307
rect 3881 23267 3939 23273
rect 5169 23307 5227 23313
rect 5169 23273 5181 23307
rect 5215 23304 5227 23307
rect 5215 23276 8064 23304
rect 5215 23273 5227 23276
rect 5169 23267 5227 23273
rect 6546 23196 6552 23248
rect 6604 23236 6610 23248
rect 6604 23208 6868 23236
rect 6604 23196 6610 23208
rect 4985 23171 5043 23177
rect 4985 23137 4997 23171
rect 5031 23168 5043 23171
rect 5258 23168 5264 23180
rect 5031 23140 5264 23168
rect 5031 23137 5043 23140
rect 4985 23131 5043 23137
rect 5258 23128 5264 23140
rect 5316 23128 5322 23180
rect 5442 23128 5448 23180
rect 5500 23168 5506 23180
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5500 23140 5825 23168
rect 5500 23128 5506 23140
rect 5813 23137 5825 23140
rect 5859 23137 5871 23171
rect 5813 23131 5871 23137
rect 5902 23128 5908 23180
rect 5960 23177 5966 23180
rect 5960 23171 6009 23177
rect 5960 23137 5963 23171
rect 5997 23137 6009 23171
rect 5960 23131 6009 23137
rect 5960 23128 5966 23131
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23168 6423 23171
rect 6638 23168 6644 23180
rect 6411 23140 6644 23168
rect 6411 23137 6423 23140
rect 6365 23131 6423 23137
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 6840 23177 6868 23208
rect 7834 23196 7840 23248
rect 7892 23196 7898 23248
rect 6825 23171 6883 23177
rect 6825 23137 6837 23171
rect 6871 23137 6883 23171
rect 6825 23131 6883 23137
rect 7006 23128 7012 23180
rect 7064 23168 7070 23180
rect 7653 23171 7711 23177
rect 7653 23168 7665 23171
rect 7064 23140 7665 23168
rect 7064 23128 7070 23140
rect 7653 23137 7665 23140
rect 7699 23137 7711 23171
rect 7653 23131 7711 23137
rect 8036 23109 8064 23276
rect 8294 23264 8300 23316
rect 8352 23264 8358 23316
rect 10045 23307 10103 23313
rect 10045 23273 10057 23307
rect 10091 23304 10103 23307
rect 12158 23304 12164 23316
rect 10091 23276 12164 23304
rect 10091 23273 10103 23276
rect 10045 23267 10103 23273
rect 12158 23264 12164 23276
rect 12216 23264 12222 23316
rect 13541 23307 13599 23313
rect 13541 23273 13553 23307
rect 13587 23304 13599 23307
rect 14734 23304 14740 23316
rect 13587 23276 14740 23304
rect 13587 23273 13599 23276
rect 13541 23267 13599 23273
rect 14734 23264 14740 23276
rect 14792 23304 14798 23316
rect 15654 23304 15660 23316
rect 14792 23276 15660 23304
rect 14792 23264 14798 23276
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16301 23307 16359 23313
rect 16301 23273 16313 23307
rect 16347 23304 16359 23307
rect 16758 23304 16764 23316
rect 16347 23276 16764 23304
rect 16347 23273 16359 23276
rect 16301 23267 16359 23273
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 17865 23307 17923 23313
rect 17865 23273 17877 23307
rect 17911 23304 17923 23307
rect 18690 23304 18696 23316
rect 17911 23276 18696 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 19886 23304 19892 23316
rect 18892 23276 19892 23304
rect 8941 23239 8999 23245
rect 8941 23205 8953 23239
rect 8987 23205 8999 23239
rect 8941 23199 8999 23205
rect 4065 23103 4123 23109
rect 4065 23069 4077 23103
rect 4111 23100 4123 23103
rect 8021 23103 8079 23109
rect 4111 23072 4384 23100
rect 4111 23069 4123 23072
rect 4065 23063 4123 23069
rect 4356 22973 4384 23072
rect 8021 23069 8033 23103
rect 8067 23069 8079 23103
rect 8021 23063 8079 23069
rect 8481 23103 8539 23109
rect 8481 23069 8493 23103
rect 8527 23100 8539 23103
rect 8956 23100 8984 23199
rect 11238 23196 11244 23248
rect 11296 23196 11302 23248
rect 11422 23196 11428 23248
rect 11480 23236 11486 23248
rect 11480 23208 11744 23236
rect 11480 23196 11486 23208
rect 9398 23128 9404 23180
rect 9456 23128 9462 23180
rect 9490 23128 9496 23180
rect 9548 23128 9554 23180
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 11716 23177 11744 23208
rect 15764 23208 15976 23236
rect 10965 23171 11023 23177
rect 10965 23168 10977 23171
rect 10100 23140 10977 23168
rect 10100 23128 10106 23140
rect 10965 23137 10977 23140
rect 11011 23137 11023 23171
rect 10965 23131 11023 23137
rect 11701 23171 11759 23177
rect 11701 23137 11713 23171
rect 11747 23137 11759 23171
rect 11701 23131 11759 23137
rect 11882 23128 11888 23180
rect 11940 23128 11946 23180
rect 15562 23128 15568 23180
rect 15620 23168 15626 23180
rect 15764 23177 15792 23208
rect 15749 23171 15807 23177
rect 15749 23168 15761 23171
rect 15620 23140 15761 23168
rect 15620 23128 15626 23140
rect 15749 23137 15761 23140
rect 15795 23137 15807 23171
rect 15749 23131 15807 23137
rect 15838 23128 15844 23180
rect 15896 23128 15902 23180
rect 15948 23168 15976 23208
rect 15948 23140 16620 23168
rect 8527 23072 8984 23100
rect 8527 23069 8539 23072
rect 8481 23063 8539 23069
rect 10686 23060 10692 23112
rect 10744 23060 10750 23112
rect 10870 23109 10876 23112
rect 10848 23103 10876 23109
rect 10848 23069 10860 23103
rect 10848 23063 10876 23069
rect 10870 23060 10876 23063
rect 10928 23060 10934 23112
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23100 12219 23103
rect 12250 23100 12256 23112
rect 12207 23072 12256 23100
rect 12207 23069 12219 23072
rect 12161 23063 12219 23069
rect 4341 22967 4399 22973
rect 4341 22933 4353 22967
rect 4387 22933 4399 22967
rect 4341 22927 4399 22933
rect 4706 22924 4712 22976
rect 4764 22924 4770 22976
rect 4798 22924 4804 22976
rect 4856 22964 4862 22976
rect 6638 22964 6644 22976
rect 4856 22936 6644 22964
rect 4856 22924 4862 22936
rect 6638 22924 6644 22936
rect 6696 22924 6702 22976
rect 6822 22924 6828 22976
rect 6880 22964 6886 22976
rect 7101 22967 7159 22973
rect 7101 22964 7113 22967
rect 6880 22936 7113 22964
rect 6880 22924 6886 22936
rect 7101 22933 7113 22936
rect 7147 22933 7159 22967
rect 7101 22927 7159 22933
rect 9309 22967 9367 22973
rect 9309 22933 9321 22967
rect 9355 22964 9367 22967
rect 9490 22964 9496 22976
rect 9355 22936 9496 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 12176 22964 12204 23063
rect 12250 23060 12256 23072
rect 12308 23060 12314 23112
rect 12434 23109 12440 23112
rect 12428 23063 12440 23109
rect 12434 23060 12440 23063
rect 12492 23060 12498 23112
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23100 14151 23103
rect 15194 23100 15200 23112
rect 14139 23072 15200 23100
rect 14139 23069 14151 23072
rect 14093 23063 14151 23069
rect 15194 23060 15200 23072
rect 15252 23100 15258 23112
rect 16206 23100 16212 23112
rect 15252 23072 16212 23100
rect 15252 23060 15258 23072
rect 16206 23060 16212 23072
rect 16264 23100 16270 23112
rect 16485 23103 16543 23109
rect 16485 23100 16497 23103
rect 16264 23072 16497 23100
rect 16264 23060 16270 23072
rect 16485 23069 16497 23072
rect 16531 23069 16543 23103
rect 16592 23100 16620 23140
rect 18414 23128 18420 23180
rect 18472 23128 18478 23180
rect 18506 23128 18512 23180
rect 18564 23128 18570 23180
rect 18230 23100 18236 23112
rect 16592 23072 18236 23100
rect 16485 23063 16543 23069
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 18322 23060 18328 23112
rect 18380 23060 18386 23112
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23100 18843 23103
rect 18892 23100 18920 23276
rect 19886 23264 19892 23276
rect 19944 23264 19950 23316
rect 19978 23264 19984 23316
rect 20036 23304 20042 23316
rect 20625 23307 20683 23313
rect 20625 23304 20637 23307
rect 20036 23276 20637 23304
rect 20036 23264 20042 23276
rect 20625 23273 20637 23276
rect 20671 23273 20683 23307
rect 20625 23267 20683 23273
rect 18831 23072 18920 23100
rect 18831 23069 18843 23072
rect 18785 23063 18843 23069
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19024 23072 19257 23100
rect 19024 23060 19030 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 14366 23041 14372 23044
rect 14360 23032 14372 23041
rect 14327 23004 14372 23032
rect 14360 22995 14372 23004
rect 14366 22992 14372 22995
rect 14424 22992 14430 23044
rect 14642 22992 14648 23044
rect 14700 23032 14706 23044
rect 15933 23035 15991 23041
rect 15933 23032 15945 23035
rect 14700 23004 15945 23032
rect 14700 22992 14706 23004
rect 15933 23001 15945 23004
rect 15979 23001 15991 23035
rect 15933 22995 15991 23001
rect 16752 23035 16810 23041
rect 16752 23001 16764 23035
rect 16798 23032 16810 23035
rect 17126 23032 17132 23044
rect 16798 23004 17132 23032
rect 16798 23001 16810 23004
rect 16752 22995 16810 23001
rect 17126 22992 17132 23004
rect 17184 22992 17190 23044
rect 17218 22992 17224 23044
rect 17276 23032 17282 23044
rect 19490 23035 19548 23041
rect 19490 23032 19502 23035
rect 17276 23004 18000 23032
rect 17276 22992 17282 23004
rect 10008 22936 12204 22964
rect 15473 22967 15531 22973
rect 10008 22924 10014 22936
rect 15473 22933 15485 22967
rect 15519 22964 15531 22967
rect 15746 22964 15752 22976
rect 15519 22936 15752 22964
rect 15519 22933 15531 22936
rect 15473 22927 15531 22933
rect 15746 22924 15752 22936
rect 15804 22964 15810 22976
rect 16390 22964 16396 22976
rect 15804 22936 16396 22964
rect 15804 22924 15810 22936
rect 16390 22924 16396 22936
rect 16448 22924 16454 22976
rect 17972 22973 18000 23004
rect 18984 23004 19502 23032
rect 18984 22973 19012 23004
rect 19490 23001 19502 23004
rect 19536 23001 19548 23035
rect 19490 22995 19548 23001
rect 17957 22967 18015 22973
rect 17957 22933 17969 22967
rect 18003 22933 18015 22967
rect 17957 22927 18015 22933
rect 18969 22967 19027 22973
rect 18969 22933 18981 22967
rect 19015 22933 19027 22967
rect 18969 22927 19027 22933
rect 1104 22874 24164 22896
rect 1104 22822 2850 22874
rect 2902 22822 2914 22874
rect 2966 22822 2978 22874
rect 3030 22822 3042 22874
rect 3094 22822 3106 22874
rect 3158 22822 5850 22874
rect 5902 22822 5914 22874
rect 5966 22822 5978 22874
rect 6030 22822 6042 22874
rect 6094 22822 6106 22874
rect 6158 22822 8850 22874
rect 8902 22822 8914 22874
rect 8966 22822 8978 22874
rect 9030 22822 9042 22874
rect 9094 22822 9106 22874
rect 9158 22822 11850 22874
rect 11902 22822 11914 22874
rect 11966 22822 11978 22874
rect 12030 22822 12042 22874
rect 12094 22822 12106 22874
rect 12158 22822 14850 22874
rect 14902 22822 14914 22874
rect 14966 22822 14978 22874
rect 15030 22822 15042 22874
rect 15094 22822 15106 22874
rect 15158 22822 17850 22874
rect 17902 22822 17914 22874
rect 17966 22822 17978 22874
rect 18030 22822 18042 22874
rect 18094 22822 18106 22874
rect 18158 22822 20850 22874
rect 20902 22822 20914 22874
rect 20966 22822 20978 22874
rect 21030 22822 21042 22874
rect 21094 22822 21106 22874
rect 21158 22822 23850 22874
rect 23902 22822 23914 22874
rect 23966 22822 23978 22874
rect 24030 22822 24042 22874
rect 24094 22822 24106 22874
rect 24158 22822 24164 22874
rect 1104 22800 24164 22822
rect 4246 22720 4252 22772
rect 4304 22720 4310 22772
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 5077 22763 5135 22769
rect 5077 22760 5089 22763
rect 4764 22732 5089 22760
rect 4764 22720 4770 22732
rect 5077 22729 5089 22732
rect 5123 22729 5135 22763
rect 5077 22723 5135 22729
rect 6270 22720 6276 22772
rect 6328 22760 6334 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 6328 22732 6377 22760
rect 6328 22720 6334 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 6365 22723 6423 22729
rect 6730 22720 6736 22772
rect 6788 22720 6794 22772
rect 6822 22720 6828 22772
rect 6880 22720 6886 22772
rect 9306 22720 9312 22772
rect 9364 22760 9370 22772
rect 9401 22763 9459 22769
rect 9401 22760 9413 22763
rect 9364 22732 9413 22760
rect 9364 22720 9370 22732
rect 9401 22729 9413 22732
rect 9447 22729 9459 22763
rect 9401 22723 9459 22729
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 10505 22763 10563 22769
rect 10505 22760 10517 22763
rect 9732 22732 10517 22760
rect 9732 22720 9738 22732
rect 10505 22729 10517 22732
rect 10551 22729 10563 22763
rect 10505 22723 10563 22729
rect 10965 22763 11023 22769
rect 10965 22729 10977 22763
rect 11011 22760 11023 22763
rect 11514 22760 11520 22772
rect 11011 22732 11520 22760
rect 11011 22729 11023 22732
rect 10965 22723 11023 22729
rect 11514 22720 11520 22732
rect 11572 22720 11578 22772
rect 13078 22720 13084 22772
rect 13136 22720 13142 22772
rect 14182 22720 14188 22772
rect 14240 22760 14246 22772
rect 14277 22763 14335 22769
rect 14277 22760 14289 22763
rect 14240 22732 14289 22760
rect 14240 22720 14246 22732
rect 14277 22729 14289 22732
rect 14323 22729 14335 22763
rect 14277 22723 14335 22729
rect 14642 22720 14648 22772
rect 14700 22720 14706 22772
rect 16850 22720 16856 22772
rect 16908 22720 16914 22772
rect 17126 22720 17132 22772
rect 17184 22720 17190 22772
rect 17586 22720 17592 22772
rect 17644 22760 17650 22772
rect 17773 22763 17831 22769
rect 17773 22760 17785 22763
rect 17644 22732 17785 22760
rect 17644 22720 17650 22732
rect 17773 22729 17785 22732
rect 17819 22729 17831 22763
rect 17773 22723 17831 22729
rect 19061 22763 19119 22769
rect 19061 22729 19073 22763
rect 19107 22760 19119 22763
rect 20254 22760 20260 22772
rect 19107 22732 20260 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 20254 22720 20260 22732
rect 20312 22720 20318 22772
rect 4617 22695 4675 22701
rect 4617 22661 4629 22695
rect 4663 22692 4675 22695
rect 4798 22692 4804 22704
rect 4663 22664 4804 22692
rect 4663 22661 4675 22664
rect 4617 22655 4675 22661
rect 4798 22652 4804 22664
rect 4856 22652 4862 22704
rect 5258 22652 5264 22704
rect 5316 22692 5322 22704
rect 8196 22695 8254 22701
rect 5316 22664 6914 22692
rect 5316 22652 5322 22664
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 4982 22624 4988 22636
rect 4755 22596 4988 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 4982 22584 4988 22596
rect 5040 22584 5046 22636
rect 5626 22584 5632 22636
rect 5684 22584 5690 22636
rect 5997 22627 6055 22633
rect 5997 22593 6009 22627
rect 6043 22624 6055 22627
rect 6362 22624 6368 22636
rect 6043 22596 6368 22624
rect 6043 22593 6055 22596
rect 5997 22587 6055 22593
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 6886 22624 6914 22664
rect 8196 22661 8208 22695
rect 8242 22692 8254 22695
rect 8386 22692 8392 22704
rect 8242 22664 8392 22692
rect 8242 22661 8254 22664
rect 8196 22655 8254 22661
rect 8386 22652 8392 22664
rect 8444 22652 8450 22704
rect 9490 22652 9496 22704
rect 9548 22692 9554 22704
rect 10873 22695 10931 22701
rect 10873 22692 10885 22695
rect 9548 22664 10885 22692
rect 9548 22652 9554 22664
rect 10873 22661 10885 22664
rect 10919 22661 10931 22695
rect 10873 22655 10931 22661
rect 13541 22695 13599 22701
rect 13541 22661 13553 22695
rect 13587 22692 13599 22695
rect 15105 22695 15163 22701
rect 15105 22692 15117 22695
rect 13587 22664 15117 22692
rect 13587 22661 13599 22664
rect 13541 22655 13599 22661
rect 15105 22661 15117 22664
rect 15151 22661 15163 22695
rect 15105 22655 15163 22661
rect 9214 22624 9220 22636
rect 6886 22596 9220 22624
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 10042 22584 10048 22636
rect 10100 22584 10106 22636
rect 13449 22627 13507 22633
rect 13449 22593 13461 22627
rect 13495 22624 13507 22627
rect 13814 22624 13820 22636
rect 13495 22596 13820 22624
rect 13495 22593 13507 22596
rect 13449 22587 13507 22593
rect 13814 22584 13820 22596
rect 13872 22624 13878 22636
rect 14642 22624 14648 22636
rect 13872 22596 14648 22624
rect 13872 22584 13878 22596
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 14737 22627 14795 22633
rect 14737 22593 14749 22627
rect 14783 22624 14795 22627
rect 15841 22627 15899 22633
rect 15841 22624 15853 22627
rect 14783 22596 15853 22624
rect 14783 22593 14795 22596
rect 14737 22587 14795 22593
rect 15841 22593 15853 22596
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 17218 22624 17224 22636
rect 17083 22596 17224 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 17310 22584 17316 22636
rect 17368 22584 17374 22636
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22624 18475 22627
rect 18690 22624 18696 22636
rect 18463 22596 18696 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 18874 22584 18880 22636
rect 18932 22584 18938 22636
rect 4890 22516 4896 22568
rect 4948 22516 4954 22568
rect 6822 22516 6828 22568
rect 6880 22556 6886 22568
rect 6917 22559 6975 22565
rect 6917 22556 6929 22559
rect 6880 22528 6929 22556
rect 6880 22516 6886 22528
rect 6917 22525 6929 22528
rect 6963 22525 6975 22559
rect 6917 22519 6975 22525
rect 7926 22516 7932 22568
rect 7984 22516 7990 22568
rect 9309 22491 9367 22497
rect 9309 22457 9321 22491
rect 9355 22488 9367 22491
rect 10060 22488 10088 22584
rect 11149 22559 11207 22565
rect 11149 22525 11161 22559
rect 11195 22525 11207 22559
rect 11149 22519 11207 22525
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22556 13783 22559
rect 14366 22556 14372 22568
rect 13771 22528 14372 22556
rect 13771 22525 13783 22528
rect 13725 22519 13783 22525
rect 9355 22460 10088 22488
rect 9355 22457 9367 22460
rect 9309 22451 9367 22457
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 5813 22423 5871 22429
rect 5813 22420 5825 22423
rect 5132 22392 5825 22420
rect 5132 22380 5138 22392
rect 5813 22389 5825 22392
rect 5859 22389 5871 22423
rect 11164 22420 11192 22519
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 14829 22559 14887 22565
rect 14829 22556 14841 22559
rect 14660 22528 14841 22556
rect 14660 22432 14688 22528
rect 14829 22525 14841 22528
rect 14875 22525 14887 22559
rect 14829 22519 14887 22525
rect 15654 22516 15660 22568
rect 15712 22516 15718 22568
rect 16390 22516 16396 22568
rect 16448 22516 16454 22568
rect 14274 22420 14280 22432
rect 11164 22392 14280 22420
rect 5813 22383 5871 22389
rect 14274 22380 14280 22392
rect 14332 22420 14338 22432
rect 14642 22420 14648 22432
rect 14332 22392 14648 22420
rect 14332 22380 14338 22392
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 1104 22330 24012 22352
rect 1104 22278 1350 22330
rect 1402 22278 1414 22330
rect 1466 22278 1478 22330
rect 1530 22278 1542 22330
rect 1594 22278 1606 22330
rect 1658 22278 4350 22330
rect 4402 22278 4414 22330
rect 4466 22278 4478 22330
rect 4530 22278 4542 22330
rect 4594 22278 4606 22330
rect 4658 22278 7350 22330
rect 7402 22278 7414 22330
rect 7466 22278 7478 22330
rect 7530 22278 7542 22330
rect 7594 22278 7606 22330
rect 7658 22278 10350 22330
rect 10402 22278 10414 22330
rect 10466 22278 10478 22330
rect 10530 22278 10542 22330
rect 10594 22278 10606 22330
rect 10658 22278 13350 22330
rect 13402 22278 13414 22330
rect 13466 22278 13478 22330
rect 13530 22278 13542 22330
rect 13594 22278 13606 22330
rect 13658 22278 16350 22330
rect 16402 22278 16414 22330
rect 16466 22278 16478 22330
rect 16530 22278 16542 22330
rect 16594 22278 16606 22330
rect 16658 22278 19350 22330
rect 19402 22278 19414 22330
rect 19466 22278 19478 22330
rect 19530 22278 19542 22330
rect 19594 22278 19606 22330
rect 19658 22278 22350 22330
rect 22402 22278 22414 22330
rect 22466 22278 22478 22330
rect 22530 22278 22542 22330
rect 22594 22278 22606 22330
rect 22658 22278 24012 22330
rect 1104 22256 24012 22278
rect 4890 22176 4896 22228
rect 4948 22216 4954 22228
rect 9398 22216 9404 22228
rect 4948 22188 9404 22216
rect 4948 22176 4954 22188
rect 5166 22040 5172 22092
rect 5224 22040 5230 22092
rect 5368 22089 5396 22188
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 9214 22108 9220 22160
rect 9272 22148 9278 22160
rect 9272 22120 9536 22148
rect 9272 22108 9278 22120
rect 5353 22083 5411 22089
rect 5353 22049 5365 22083
rect 5399 22049 5411 22083
rect 5353 22043 5411 22049
rect 6917 22083 6975 22089
rect 6917 22049 6929 22083
rect 6963 22080 6975 22083
rect 7926 22080 7932 22092
rect 6963 22052 7932 22080
rect 6963 22049 6975 22052
rect 6917 22043 6975 22049
rect 4614 21972 4620 22024
rect 4672 21972 4678 22024
rect 4798 21904 4804 21956
rect 4856 21944 4862 21956
rect 5077 21947 5135 21953
rect 5077 21944 5089 21947
rect 4856 21916 5089 21944
rect 4856 21904 4862 21916
rect 5077 21913 5089 21916
rect 5123 21944 5135 21947
rect 5184 21944 5212 22040
rect 5626 21972 5632 22024
rect 5684 22012 5690 22024
rect 6089 22015 6147 22021
rect 6089 22012 6101 22015
rect 5684 21984 6101 22012
rect 5684 21972 5690 21984
rect 6089 21981 6101 21984
rect 6135 21981 6147 22015
rect 6089 21975 6147 21981
rect 6549 22015 6607 22021
rect 6549 21981 6561 22015
rect 6595 22012 6607 22015
rect 6932 22012 6960 22043
rect 7926 22040 7932 22052
rect 7984 22040 7990 22092
rect 9508 22089 9536 22120
rect 13722 22108 13728 22160
rect 13780 22148 13786 22160
rect 18414 22148 18420 22160
rect 13780 22120 18420 22148
rect 13780 22108 13786 22120
rect 18414 22108 18420 22120
rect 18472 22108 18478 22160
rect 9493 22083 9551 22089
rect 9493 22080 9505 22083
rect 9471 22052 9505 22080
rect 9493 22049 9505 22052
rect 9539 22049 9551 22083
rect 9493 22043 9551 22049
rect 14182 22040 14188 22092
rect 14240 22080 14246 22092
rect 14366 22080 14372 22092
rect 14240 22052 14372 22080
rect 14240 22040 14246 22052
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 6595 21984 6960 22012
rect 6595 21981 6607 21984
rect 6549 21975 6607 21981
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 9398 22012 9404 22024
rect 8812 21984 9404 22012
rect 8812 21972 8818 21984
rect 9398 21972 9404 21984
rect 9456 21972 9462 22024
rect 10318 21972 10324 22024
rect 10376 21972 10382 22024
rect 10689 22015 10747 22021
rect 10689 21981 10701 22015
rect 10735 22012 10747 22015
rect 11514 22012 11520 22024
rect 10735 21984 11520 22012
rect 10735 21981 10747 21984
rect 10689 21975 10747 21981
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 22012 12955 22015
rect 13170 22012 13176 22024
rect 12943 21984 13176 22012
rect 12943 21981 12955 21984
rect 12897 21975 12955 21981
rect 6730 21944 6736 21956
rect 5123 21916 6736 21944
rect 5123 21913 5135 21916
rect 5077 21907 5135 21913
rect 6730 21904 6736 21916
rect 6788 21904 6794 21956
rect 7650 21904 7656 21956
rect 7708 21904 7714 21956
rect 9309 21947 9367 21953
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 9769 21947 9827 21953
rect 9769 21944 9781 21947
rect 9355 21916 9781 21944
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 9769 21913 9781 21916
rect 9815 21913 9827 21947
rect 12636 21944 12664 21975
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 14734 21972 14740 22024
rect 14792 21972 14798 22024
rect 15378 21972 15384 22024
rect 15436 21972 15442 22024
rect 16666 21972 16672 22024
rect 16724 21972 16730 22024
rect 19061 22015 19119 22021
rect 19061 21981 19073 22015
rect 19107 22012 19119 22015
rect 19242 22012 19248 22024
rect 19107 21984 19248 22012
rect 19107 21981 19119 21984
rect 19061 21975 19119 21981
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 13998 21944 14004 21956
rect 12636 21916 14004 21944
rect 9769 21907 9827 21913
rect 13998 21904 14004 21916
rect 14056 21904 14062 21956
rect 16298 21904 16304 21956
rect 16356 21944 16362 21956
rect 18966 21944 18972 21956
rect 16356 21916 18972 21944
rect 16356 21904 16362 21916
rect 18966 21904 18972 21916
rect 19024 21904 19030 21956
rect 3973 21879 4031 21885
rect 3973 21845 3985 21879
rect 4019 21876 4031 21879
rect 4246 21876 4252 21888
rect 4019 21848 4252 21876
rect 4019 21845 4031 21848
rect 3973 21839 4031 21845
rect 4246 21836 4252 21848
rect 4304 21836 4310 21888
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 5169 21879 5227 21885
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5537 21879 5595 21885
rect 5537 21876 5549 21879
rect 5215 21848 5549 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5537 21845 5549 21848
rect 5583 21845 5595 21879
rect 5537 21839 5595 21845
rect 7929 21879 7987 21885
rect 7929 21845 7941 21879
rect 7975 21876 7987 21879
rect 8018 21876 8024 21888
rect 7975 21848 8024 21876
rect 7975 21845 7987 21848
rect 7929 21839 7987 21845
rect 8018 21836 8024 21848
rect 8076 21836 8082 21888
rect 8941 21879 8999 21885
rect 8941 21845 8953 21879
rect 8987 21876 8999 21879
rect 9214 21876 9220 21888
rect 8987 21848 9220 21876
rect 8987 21845 8999 21848
rect 8941 21839 8999 21845
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 10226 21836 10232 21888
rect 10284 21876 10290 21888
rect 10505 21879 10563 21885
rect 10505 21876 10517 21879
rect 10284 21848 10517 21876
rect 10284 21836 10290 21848
rect 10505 21845 10517 21848
rect 10551 21845 10563 21879
rect 10505 21839 10563 21845
rect 12437 21879 12495 21885
rect 12437 21845 12449 21879
rect 12483 21876 12495 21879
rect 12526 21876 12532 21888
rect 12483 21848 12532 21876
rect 12483 21845 12495 21848
rect 12437 21839 12495 21845
rect 12526 21836 12532 21848
rect 12584 21836 12590 21888
rect 12710 21836 12716 21888
rect 12768 21836 12774 21888
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 13596 21848 14105 21876
rect 13596 21836 13602 21848
rect 14093 21845 14105 21848
rect 14139 21845 14151 21879
rect 14093 21839 14151 21845
rect 14458 21836 14464 21888
rect 14516 21876 14522 21888
rect 14829 21879 14887 21885
rect 14829 21876 14841 21879
rect 14516 21848 14841 21876
rect 14516 21836 14522 21848
rect 14829 21845 14841 21848
rect 14875 21845 14887 21879
rect 14829 21839 14887 21845
rect 15654 21836 15660 21888
rect 15712 21876 15718 21888
rect 16117 21879 16175 21885
rect 16117 21876 16129 21879
rect 15712 21848 16129 21876
rect 15712 21836 15718 21848
rect 16117 21845 16129 21848
rect 16163 21845 16175 21879
rect 16117 21839 16175 21845
rect 18417 21879 18475 21885
rect 18417 21845 18429 21879
rect 18463 21876 18475 21879
rect 18506 21876 18512 21888
rect 18463 21848 18512 21876
rect 18463 21845 18475 21848
rect 18417 21839 18475 21845
rect 18506 21836 18512 21848
rect 18564 21836 18570 21888
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 19705 21879 19763 21885
rect 19705 21876 19717 21879
rect 18656 21848 19717 21876
rect 18656 21836 18662 21848
rect 19705 21845 19717 21848
rect 19751 21845 19763 21879
rect 19705 21839 19763 21845
rect 1104 21786 24164 21808
rect 1104 21734 2850 21786
rect 2902 21734 2914 21786
rect 2966 21734 2978 21786
rect 3030 21734 3042 21786
rect 3094 21734 3106 21786
rect 3158 21734 5850 21786
rect 5902 21734 5914 21786
rect 5966 21734 5978 21786
rect 6030 21734 6042 21786
rect 6094 21734 6106 21786
rect 6158 21734 8850 21786
rect 8902 21734 8914 21786
rect 8966 21734 8978 21786
rect 9030 21734 9042 21786
rect 9094 21734 9106 21786
rect 9158 21734 11850 21786
rect 11902 21734 11914 21786
rect 11966 21734 11978 21786
rect 12030 21734 12042 21786
rect 12094 21734 12106 21786
rect 12158 21734 14850 21786
rect 14902 21734 14914 21786
rect 14966 21734 14978 21786
rect 15030 21734 15042 21786
rect 15094 21734 15106 21786
rect 15158 21734 17850 21786
rect 17902 21734 17914 21786
rect 17966 21734 17978 21786
rect 18030 21734 18042 21786
rect 18094 21734 18106 21786
rect 18158 21734 20850 21786
rect 20902 21734 20914 21786
rect 20966 21734 20978 21786
rect 21030 21734 21042 21786
rect 21094 21734 21106 21786
rect 21158 21734 23850 21786
rect 23902 21734 23914 21786
rect 23966 21734 23978 21786
rect 24030 21734 24042 21786
rect 24094 21734 24106 21786
rect 24158 21734 24164 21786
rect 1104 21712 24164 21734
rect 6362 21632 6368 21684
rect 6420 21632 6426 21684
rect 11514 21632 11520 21684
rect 11572 21632 11578 21684
rect 13170 21632 13176 21684
rect 13228 21632 13234 21684
rect 13538 21632 13544 21684
rect 13596 21632 13602 21684
rect 13998 21632 14004 21684
rect 14056 21632 14062 21684
rect 14458 21632 14464 21684
rect 14516 21632 14522 21684
rect 14642 21632 14648 21684
rect 14700 21672 14706 21684
rect 15013 21675 15071 21681
rect 15013 21672 15025 21675
rect 14700 21644 15025 21672
rect 14700 21632 14706 21644
rect 15013 21641 15025 21644
rect 15059 21672 15071 21675
rect 16666 21672 16672 21684
rect 15059 21644 16672 21672
rect 15059 21641 15071 21644
rect 15013 21635 15071 21641
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 17678 21672 17684 21684
rect 16776 21644 17684 21672
rect 5166 21564 5172 21616
rect 5224 21564 5230 21616
rect 9398 21564 9404 21616
rect 9456 21604 9462 21616
rect 11885 21607 11943 21613
rect 11885 21604 11897 21607
rect 9456 21576 11897 21604
rect 9456 21564 9462 21576
rect 11885 21573 11897 21576
rect 11931 21573 11943 21607
rect 16776 21604 16804 21644
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 18598 21632 18604 21684
rect 18656 21632 18662 21684
rect 18690 21632 18696 21684
rect 18748 21672 18754 21684
rect 20438 21672 20444 21684
rect 18748 21644 20444 21672
rect 18748 21632 18754 21644
rect 20438 21632 20444 21644
rect 20496 21632 20502 21684
rect 11885 21567 11943 21573
rect 15396 21576 16804 21604
rect 3504 21539 3562 21545
rect 3504 21505 3516 21539
rect 3550 21536 3562 21539
rect 3786 21536 3792 21548
rect 3550 21508 3792 21536
rect 3550 21505 3562 21508
rect 3504 21499 3562 21505
rect 3786 21496 3792 21508
rect 3844 21496 3850 21548
rect 5077 21539 5135 21545
rect 5077 21505 5089 21539
rect 5123 21505 5135 21539
rect 5077 21499 5135 21505
rect 3237 21471 3295 21477
rect 3237 21437 3249 21471
rect 3283 21437 3295 21471
rect 5092 21468 5120 21499
rect 6730 21496 6736 21548
rect 6788 21496 6794 21548
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21536 6883 21539
rect 7193 21539 7251 21545
rect 7193 21536 7205 21539
rect 6871 21508 7205 21536
rect 6871 21505 6883 21508
rect 6825 21499 6883 21505
rect 7193 21505 7205 21508
rect 7239 21505 7251 21539
rect 7193 21499 7251 21505
rect 8288 21539 8346 21545
rect 8288 21505 8300 21539
rect 8334 21536 8346 21539
rect 8846 21536 8852 21548
rect 8334 21508 8852 21536
rect 8334 21505 8346 21508
rect 8288 21499 8346 21505
rect 8846 21496 8852 21508
rect 8904 21496 8910 21548
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10209 21539 10267 21545
rect 10209 21536 10221 21539
rect 10060 21508 10221 21536
rect 5442 21468 5448 21480
rect 5092 21440 5448 21468
rect 3237 21431 3295 21437
rect 3252 21332 3280 21431
rect 5442 21428 5448 21440
rect 5500 21468 5506 21480
rect 5905 21471 5963 21477
rect 5905 21468 5917 21471
rect 5500 21440 5917 21468
rect 5500 21428 5506 21440
rect 5905 21437 5917 21440
rect 5951 21437 5963 21471
rect 5905 21431 5963 21437
rect 6638 21428 6644 21480
rect 6696 21468 6702 21480
rect 6917 21471 6975 21477
rect 6917 21468 6929 21471
rect 6696 21440 6929 21468
rect 6696 21428 6702 21440
rect 6917 21437 6929 21440
rect 6963 21437 6975 21471
rect 6917 21431 6975 21437
rect 7006 21428 7012 21480
rect 7064 21468 7070 21480
rect 7745 21471 7803 21477
rect 7745 21468 7757 21471
rect 7064 21440 7757 21468
rect 7064 21428 7070 21440
rect 7745 21437 7757 21440
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 7926 21428 7932 21480
rect 7984 21468 7990 21480
rect 8021 21471 8079 21477
rect 8021 21468 8033 21471
rect 7984 21440 8033 21468
rect 7984 21428 7990 21440
rect 8021 21437 8033 21440
rect 8067 21437 8079 21471
rect 8021 21431 8079 21437
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10060 21468 10088 21508
rect 10209 21505 10221 21508
rect 10255 21505 10267 21539
rect 10209 21499 10267 21505
rect 11977 21539 12035 21545
rect 11977 21505 11989 21539
rect 12023 21536 12035 21539
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 12023 21508 12357 21536
rect 12023 21505 12035 21508
rect 11977 21499 12035 21505
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 13633 21539 13691 21545
rect 13633 21505 13645 21539
rect 13679 21536 13691 21539
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 13679 21508 14381 21536
rect 13679 21505 13691 21508
rect 13633 21499 13691 21505
rect 14369 21505 14381 21508
rect 14415 21536 14427 21539
rect 14458 21536 14464 21548
rect 14415 21508 14464 21536
rect 14415 21505 14427 21508
rect 14369 21499 14427 21505
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 9732 21440 10088 21468
rect 9732 21428 9738 21440
rect 11514 21428 11520 21480
rect 11572 21468 11578 21480
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 11572 21440 12081 21468
rect 11572 21428 11578 21440
rect 12069 21437 12081 21440
rect 12115 21437 12127 21471
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12069 21431 12127 21437
rect 12406 21440 12909 21468
rect 11422 21360 11428 21412
rect 11480 21400 11486 21412
rect 12406 21400 12434 21440
rect 12897 21437 12909 21440
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 13722 21428 13728 21480
rect 13780 21428 13786 21480
rect 14182 21428 14188 21480
rect 14240 21468 14246 21480
rect 14645 21471 14703 21477
rect 14645 21468 14657 21471
rect 14240 21440 14657 21468
rect 14240 21428 14246 21440
rect 14645 21437 14657 21440
rect 14691 21468 14703 21471
rect 15396 21468 15424 21576
rect 16114 21496 16120 21548
rect 16172 21545 16178 21548
rect 16172 21499 16184 21545
rect 16172 21496 16178 21499
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 16393 21539 16451 21545
rect 16393 21536 16405 21539
rect 16356 21508 16405 21536
rect 16356 21496 16362 21508
rect 16393 21505 16405 21508
rect 16439 21536 16451 21539
rect 16761 21539 16819 21545
rect 16761 21536 16773 21539
rect 16439 21508 16773 21536
rect 16439 21505 16451 21508
rect 16393 21499 16451 21505
rect 16761 21505 16773 21508
rect 16807 21505 16819 21539
rect 16761 21499 16819 21505
rect 16850 21496 16856 21548
rect 16908 21536 16914 21548
rect 17017 21539 17075 21545
rect 17017 21536 17029 21539
rect 16908 21508 17029 21536
rect 16908 21496 16914 21508
rect 17017 21505 17029 21508
rect 17063 21505 17075 21539
rect 17017 21499 17075 21505
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 18782 21536 18788 21548
rect 18739 21508 18788 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 18966 21496 18972 21548
rect 19024 21536 19030 21548
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 19024 21508 19165 21536
rect 19024 21496 19030 21508
rect 19153 21505 19165 21508
rect 19199 21505 19211 21539
rect 19153 21499 19211 21505
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 19420 21539 19478 21545
rect 19420 21505 19432 21539
rect 19466 21536 19478 21539
rect 19978 21536 19984 21548
rect 19466 21508 19984 21536
rect 19466 21505 19478 21508
rect 19420 21499 19478 21505
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 21324 21508 23397 21536
rect 21324 21496 21330 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 18417 21471 18475 21477
rect 18417 21468 18429 21471
rect 14691 21440 15424 21468
rect 17880 21440 18429 21468
rect 14691 21437 14703 21440
rect 14645 21431 14703 21437
rect 11480 21372 12434 21400
rect 11480 21360 11486 21372
rect 4154 21332 4160 21344
rect 3252 21304 4160 21332
rect 4154 21292 4160 21304
rect 4212 21292 4218 21344
rect 4614 21292 4620 21344
rect 4672 21332 4678 21344
rect 6086 21332 6092 21344
rect 4672 21304 6092 21332
rect 4672 21292 4678 21304
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 9401 21335 9459 21341
rect 9401 21301 9413 21335
rect 9447 21332 9459 21335
rect 10134 21332 10140 21344
rect 9447 21304 10140 21332
rect 9447 21301 9459 21304
rect 9401 21295 9459 21301
rect 10134 21292 10140 21304
rect 10192 21332 10198 21344
rect 10318 21332 10324 21344
rect 10192 21304 10324 21332
rect 10192 21292 10198 21304
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 11330 21292 11336 21344
rect 11388 21292 11394 21344
rect 14550 21292 14556 21344
rect 14608 21332 14614 21344
rect 17880 21332 17908 21440
rect 18417 21437 18429 21440
rect 18463 21468 18475 21471
rect 18598 21468 18604 21480
rect 18463 21440 18604 21468
rect 18463 21437 18475 21440
rect 18417 21431 18475 21437
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 19260 21468 19288 21496
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 18708 21440 19288 21468
rect 20548 21440 20913 21468
rect 18141 21403 18199 21409
rect 18141 21369 18153 21403
rect 18187 21400 18199 21403
rect 18708 21400 18736 21440
rect 18187 21372 18736 21400
rect 18187 21369 18199 21372
rect 18141 21363 18199 21369
rect 14608 21304 17908 21332
rect 19061 21335 19119 21341
rect 14608 21292 14614 21304
rect 19061 21301 19073 21335
rect 19107 21332 19119 21335
rect 19150 21332 19156 21344
rect 19107 21304 19156 21332
rect 19107 21301 19119 21304
rect 19061 21295 19119 21301
rect 19150 21292 19156 21304
rect 19208 21292 19214 21344
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 20548 21341 20576 21440
rect 20901 21437 20913 21440
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 20533 21335 20591 21341
rect 20533 21332 20545 21335
rect 19852 21304 20545 21332
rect 19852 21292 19858 21304
rect 20533 21301 20545 21304
rect 20579 21301 20591 21335
rect 20533 21295 20591 21301
rect 21174 21292 21180 21344
rect 21232 21332 21238 21344
rect 21545 21335 21603 21341
rect 21545 21332 21557 21335
rect 21232 21304 21557 21332
rect 21232 21292 21238 21304
rect 21545 21301 21557 21304
rect 21591 21301 21603 21335
rect 21545 21295 21603 21301
rect 23566 21292 23572 21344
rect 23624 21292 23630 21344
rect 1104 21242 24012 21264
rect 1104 21190 1350 21242
rect 1402 21190 1414 21242
rect 1466 21190 1478 21242
rect 1530 21190 1542 21242
rect 1594 21190 1606 21242
rect 1658 21190 4350 21242
rect 4402 21190 4414 21242
rect 4466 21190 4478 21242
rect 4530 21190 4542 21242
rect 4594 21190 4606 21242
rect 4658 21190 7350 21242
rect 7402 21190 7414 21242
rect 7466 21190 7478 21242
rect 7530 21190 7542 21242
rect 7594 21190 7606 21242
rect 7658 21190 10350 21242
rect 10402 21190 10414 21242
rect 10466 21190 10478 21242
rect 10530 21190 10542 21242
rect 10594 21190 10606 21242
rect 10658 21190 13350 21242
rect 13402 21190 13414 21242
rect 13466 21190 13478 21242
rect 13530 21190 13542 21242
rect 13594 21190 13606 21242
rect 13658 21190 16350 21242
rect 16402 21190 16414 21242
rect 16466 21190 16478 21242
rect 16530 21190 16542 21242
rect 16594 21190 16606 21242
rect 16658 21190 19350 21242
rect 19402 21190 19414 21242
rect 19466 21190 19478 21242
rect 19530 21190 19542 21242
rect 19594 21190 19606 21242
rect 19658 21190 22350 21242
rect 22402 21190 22414 21242
rect 22466 21190 22478 21242
rect 22530 21190 22542 21242
rect 22594 21190 22606 21242
rect 22658 21190 24012 21242
rect 1104 21168 24012 21190
rect 3786 21088 3792 21140
rect 3844 21088 3850 21140
rect 4706 21128 4712 21140
rect 4632 21100 4712 21128
rect 4632 21060 4660 21100
rect 4706 21088 4712 21100
rect 4764 21088 4770 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8904 21100 8953 21128
rect 8904 21088 8910 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 10134 21088 10140 21140
rect 10192 21128 10198 21140
rect 10192 21100 10456 21128
rect 10192 21088 10198 21100
rect 3620 21032 4660 21060
rect 3620 20933 3648 21032
rect 6546 21020 6552 21072
rect 6604 21020 6610 21072
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20992 4767 20995
rect 5258 20992 5264 21004
rect 4755 20964 5264 20992
rect 4755 20961 4767 20964
rect 4709 20955 4767 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 5951 20995 6009 21001
rect 5951 20992 5963 20995
rect 5684 20964 5963 20992
rect 5684 20952 5690 20964
rect 5951 20961 5963 20964
rect 5997 20961 6009 20995
rect 5951 20955 6009 20961
rect 6086 20952 6092 21004
rect 6144 20952 6150 21004
rect 6270 20952 6276 21004
rect 6328 20992 6334 21004
rect 6365 20995 6423 21001
rect 6365 20992 6377 20995
rect 6328 20964 6377 20992
rect 6328 20952 6334 20964
rect 6365 20961 6377 20964
rect 6411 20992 6423 20995
rect 6564 20992 6592 21020
rect 6411 20964 6592 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 7006 20952 7012 21004
rect 7064 20952 7070 21004
rect 9306 20952 9312 21004
rect 9364 20992 9370 21004
rect 10112 20995 10170 21001
rect 10112 20992 10124 20995
rect 9364 20964 10124 20992
rect 9364 20952 9370 20964
rect 10112 20961 10124 20964
rect 10158 20961 10170 20995
rect 10428 20992 10456 21100
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 14148 21100 14734 21128
rect 14148 21088 14154 21100
rect 13630 21020 13636 21072
rect 13688 21020 13694 21072
rect 14550 21060 14556 21072
rect 14292 21032 14556 21060
rect 10112 20955 10170 20961
rect 10244 20964 10456 20992
rect 10505 20995 10563 21001
rect 3605 20927 3663 20933
rect 3605 20893 3617 20927
rect 3651 20893 3663 20927
rect 3605 20887 3663 20893
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20924 4031 20927
rect 4019 20896 4200 20924
rect 4019 20893 4031 20896
rect 3973 20887 4031 20893
rect 3421 20791 3479 20797
rect 3421 20757 3433 20791
rect 3467 20788 3479 20791
rect 3510 20788 3516 20800
rect 3467 20760 3516 20788
rect 3467 20757 3479 20760
rect 3421 20751 3479 20757
rect 3510 20748 3516 20760
rect 3568 20748 3574 20800
rect 4172 20797 4200 20896
rect 4246 20884 4252 20936
rect 4304 20924 4310 20936
rect 4525 20927 4583 20933
rect 4525 20924 4537 20927
rect 4304 20896 4537 20924
rect 4304 20884 4310 20896
rect 4525 20893 4537 20896
rect 4571 20893 4583 20927
rect 4525 20887 4583 20893
rect 4617 20927 4675 20933
rect 4617 20893 4629 20927
rect 4663 20924 4675 20927
rect 4798 20924 4804 20936
rect 4663 20896 4804 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 4157 20791 4215 20797
rect 4157 20757 4169 20791
rect 4203 20757 4215 20791
rect 4157 20751 4215 20757
rect 5169 20791 5227 20797
rect 5169 20757 5181 20791
rect 5215 20788 5227 20791
rect 6638 20788 6644 20800
rect 5215 20760 6644 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 6840 20788 6868 20887
rect 7926 20884 7932 20936
rect 7984 20924 7990 20936
rect 8481 20927 8539 20933
rect 8481 20924 8493 20927
rect 7984 20896 8493 20924
rect 7984 20884 7990 20896
rect 8481 20893 8493 20896
rect 8527 20893 8539 20927
rect 8481 20887 8539 20893
rect 8754 20884 8760 20936
rect 8812 20884 8818 20936
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20924 9183 20927
rect 9214 20924 9220 20936
rect 9171 20896 9220 20924
rect 9171 20893 9183 20896
rect 9125 20887 9183 20893
rect 9214 20884 9220 20896
rect 9272 20884 9278 20936
rect 9950 20884 9956 20936
rect 10008 20884 10014 20936
rect 10244 20933 10272 20964
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 10870 20992 10876 21004
rect 10551 20964 10876 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 10870 20952 10876 20964
rect 10928 20952 10934 21004
rect 10965 20995 11023 21001
rect 10965 20961 10977 20995
rect 11011 20992 11023 20995
rect 11330 20992 11336 21004
rect 11011 20964 11336 20992
rect 11011 20961 11023 20964
rect 10965 20955 11023 20961
rect 11330 20952 11336 20964
rect 11388 20952 11394 21004
rect 14292 21001 14320 21032
rect 14550 21020 14556 21032
rect 14608 21020 14614 21072
rect 14706 21001 14734 21100
rect 15102 21088 15108 21140
rect 15160 21128 15166 21140
rect 15378 21128 15384 21140
rect 15160 21100 15384 21128
rect 15160 21088 15166 21100
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16209 21131 16267 21137
rect 16209 21128 16221 21131
rect 16080 21100 16221 21128
rect 16080 21088 16086 21100
rect 16209 21097 16221 21100
rect 16255 21097 16267 21131
rect 16209 21091 16267 21097
rect 16577 21131 16635 21137
rect 16577 21097 16589 21131
rect 16623 21128 16635 21131
rect 16850 21128 16856 21140
rect 16623 21100 16856 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 20346 21088 20352 21140
rect 20404 21128 20410 21140
rect 20625 21131 20683 21137
rect 20625 21128 20637 21131
rect 20404 21100 20637 21128
rect 20404 21088 20410 21100
rect 20625 21097 20637 21100
rect 20671 21097 20683 21131
rect 20625 21091 20683 21097
rect 18049 21063 18107 21069
rect 18049 21029 18061 21063
rect 18095 21060 18107 21063
rect 18966 21060 18972 21072
rect 18095 21032 18972 21060
rect 18095 21029 18107 21032
rect 18049 21023 18107 21029
rect 18966 21020 18972 21032
rect 19024 21020 19030 21072
rect 14277 20995 14335 21001
rect 14277 20961 14289 20995
rect 14323 20961 14335 20995
rect 14706 20995 14775 21001
rect 14706 20964 14729 20995
rect 14277 20955 14335 20961
rect 14717 20961 14729 20964
rect 14763 20961 14775 20995
rect 14717 20955 14775 20961
rect 15102 20952 15108 21004
rect 15160 21001 15166 21004
rect 15160 20995 15188 21001
rect 15176 20961 15188 20995
rect 15160 20955 15188 20961
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20992 15347 20995
rect 15470 20992 15476 21004
rect 15335 20964 15476 20992
rect 15335 20961 15347 20964
rect 15289 20955 15347 20961
rect 15160 20952 15166 20955
rect 15470 20952 15476 20964
rect 15528 20992 15534 21004
rect 15838 20992 15844 21004
rect 15528 20964 15844 20992
rect 15528 20952 15534 20964
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 18414 20952 18420 21004
rect 18472 20992 18478 21004
rect 18693 20995 18751 21001
rect 18693 20992 18705 20995
rect 18472 20964 18705 20992
rect 18472 20952 18478 20964
rect 18693 20961 18705 20964
rect 18739 20961 18751 20995
rect 18693 20955 18751 20961
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 19116 20964 19257 20992
rect 19116 20952 19122 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 19245 20955 19303 20961
rect 21174 20952 21180 21004
rect 21232 20952 21238 21004
rect 21358 20952 21364 21004
rect 21416 20952 21422 21004
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20893 11207 20927
rect 11149 20887 11207 20893
rect 8018 20816 8024 20868
rect 8076 20856 8082 20868
rect 8214 20859 8272 20865
rect 8214 20856 8226 20859
rect 8076 20828 8226 20856
rect 8076 20816 8082 20828
rect 8214 20825 8226 20828
rect 8260 20825 8272 20859
rect 11164 20856 11192 20887
rect 11238 20884 11244 20936
rect 11296 20884 11302 20936
rect 12526 20933 12532 20936
rect 12242 20927 12300 20933
rect 12242 20924 12254 20927
rect 11992 20896 12254 20924
rect 11422 20856 11428 20868
rect 11164 20828 11428 20856
rect 8214 20819 8272 20825
rect 11422 20816 11428 20828
rect 11480 20816 11486 20868
rect 11992 20865 12020 20896
rect 12242 20893 12254 20896
rect 12288 20893 12300 20927
rect 12242 20887 12300 20893
rect 12520 20887 12532 20933
rect 12526 20884 12532 20887
rect 12584 20884 12590 20936
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 13906 20924 13912 20936
rect 13771 20896 13912 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 13906 20884 13912 20896
rect 13964 20884 13970 20936
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 11977 20859 12035 20865
rect 11977 20825 11989 20859
rect 12023 20825 12035 20859
rect 11977 20819 12035 20825
rect 7098 20788 7104 20800
rect 6840 20760 7104 20788
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 8570 20748 8576 20800
rect 8628 20748 8634 20800
rect 9309 20791 9367 20797
rect 9309 20757 9321 20791
rect 9355 20788 9367 20791
rect 11146 20788 11152 20800
rect 9355 20760 11152 20788
rect 9355 20757 9367 20760
rect 9309 20751 9367 20757
rect 11146 20748 11152 20760
rect 11204 20748 11210 20800
rect 11238 20748 11244 20800
rect 11296 20788 11302 20800
rect 11992 20788 12020 20819
rect 11296 20760 12020 20788
rect 13909 20791 13967 20797
rect 11296 20748 11302 20760
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 13998 20788 14004 20800
rect 13955 20760 14004 20788
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 13998 20748 14004 20760
rect 14056 20748 14062 20800
rect 14108 20788 14136 20887
rect 15010 20884 15016 20936
rect 15068 20884 15074 20936
rect 15933 20927 15991 20933
rect 15933 20893 15945 20927
rect 15979 20924 15991 20927
rect 16025 20927 16083 20933
rect 16025 20924 16037 20927
rect 15979 20896 16037 20924
rect 15979 20893 15991 20896
rect 15933 20887 15991 20893
rect 16025 20893 16037 20896
rect 16071 20893 16083 20927
rect 16025 20887 16083 20893
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 16408 20856 16436 20887
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 16669 20927 16727 20933
rect 16669 20924 16681 20927
rect 16540 20896 16681 20924
rect 16540 20884 16546 20896
rect 16669 20893 16681 20896
rect 16715 20893 16727 20927
rect 16669 20887 16727 20893
rect 16776 20896 18184 20924
rect 16776 20856 16804 20896
rect 16942 20865 16948 20868
rect 16408 20828 16804 20856
rect 16936 20819 16948 20865
rect 16942 20816 16948 20819
rect 17000 20816 17006 20868
rect 15378 20788 15384 20800
rect 14108 20760 15384 20788
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 18156 20797 18184 20896
rect 18506 20884 18512 20936
rect 18564 20884 18570 20936
rect 20714 20884 20720 20936
rect 20772 20884 20778 20936
rect 19512 20859 19570 20865
rect 19512 20825 19524 20859
rect 19558 20856 19570 20859
rect 19702 20856 19708 20868
rect 19558 20828 19708 20856
rect 19558 20825 19570 20828
rect 19512 20819 19570 20825
rect 19702 20816 19708 20828
rect 19760 20816 19766 20868
rect 20732 20856 20760 20884
rect 21085 20859 21143 20865
rect 21085 20856 21097 20859
rect 19812 20828 21097 20856
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20757 18199 20791
rect 18141 20751 18199 20757
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 19812 20788 19840 20828
rect 21085 20825 21097 20828
rect 21131 20825 21143 20859
rect 21085 20819 21143 20825
rect 18656 20760 19840 20788
rect 18656 20748 18662 20760
rect 20714 20748 20720 20800
rect 20772 20748 20778 20800
rect 1104 20698 24164 20720
rect 1104 20646 2850 20698
rect 2902 20646 2914 20698
rect 2966 20646 2978 20698
rect 3030 20646 3042 20698
rect 3094 20646 3106 20698
rect 3158 20646 5850 20698
rect 5902 20646 5914 20698
rect 5966 20646 5978 20698
rect 6030 20646 6042 20698
rect 6094 20646 6106 20698
rect 6158 20646 8850 20698
rect 8902 20646 8914 20698
rect 8966 20646 8978 20698
rect 9030 20646 9042 20698
rect 9094 20646 9106 20698
rect 9158 20646 11850 20698
rect 11902 20646 11914 20698
rect 11966 20646 11978 20698
rect 12030 20646 12042 20698
rect 12094 20646 12106 20698
rect 12158 20646 14850 20698
rect 14902 20646 14914 20698
rect 14966 20646 14978 20698
rect 15030 20646 15042 20698
rect 15094 20646 15106 20698
rect 15158 20646 17850 20698
rect 17902 20646 17914 20698
rect 17966 20646 17978 20698
rect 18030 20646 18042 20698
rect 18094 20646 18106 20698
rect 18158 20646 20850 20698
rect 20902 20646 20914 20698
rect 20966 20646 20978 20698
rect 21030 20646 21042 20698
rect 21094 20646 21106 20698
rect 21158 20646 23850 20698
rect 23902 20646 23914 20698
rect 23966 20646 23978 20698
rect 24030 20646 24042 20698
rect 24094 20646 24106 20698
rect 24158 20646 24164 20698
rect 1104 20624 24164 20646
rect 4617 20587 4675 20593
rect 4617 20553 4629 20587
rect 4663 20584 4675 20587
rect 5626 20584 5632 20596
rect 4663 20556 5632 20584
rect 4663 20553 4675 20556
rect 4617 20547 4675 20553
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 6181 20587 6239 20593
rect 6181 20553 6193 20587
rect 6227 20584 6239 20587
rect 7006 20584 7012 20596
rect 6227 20556 7012 20584
rect 6227 20553 6239 20556
rect 6181 20547 6239 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 7101 20587 7159 20593
rect 7101 20553 7113 20587
rect 7147 20584 7159 20587
rect 7742 20584 7748 20596
rect 7147 20556 7748 20584
rect 7147 20553 7159 20556
rect 7101 20547 7159 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 9306 20544 9312 20596
rect 9364 20544 9370 20596
rect 9861 20587 9919 20593
rect 9861 20553 9873 20587
rect 9907 20553 9919 20587
rect 9861 20547 9919 20553
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 11422 20584 11428 20596
rect 11379 20556 11428 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 5442 20516 5448 20528
rect 4816 20488 5448 20516
rect 3510 20457 3516 20460
rect 3504 20448 3516 20457
rect 3471 20420 3516 20448
rect 3504 20411 3516 20420
rect 3510 20408 3516 20411
rect 3568 20408 3574 20460
rect 4816 20389 4844 20488
rect 5442 20476 5448 20488
rect 5500 20516 5506 20528
rect 8196 20519 8254 20525
rect 5500 20488 7972 20516
rect 5500 20476 5506 20488
rect 5074 20457 5080 20460
rect 5068 20448 5080 20457
rect 5035 20420 5080 20448
rect 5068 20411 5080 20420
rect 5074 20408 5080 20411
rect 5132 20408 5138 20460
rect 6730 20408 6736 20460
rect 6788 20408 6794 20460
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7944 20457 7972 20488
rect 8196 20485 8208 20519
rect 8242 20516 8254 20519
rect 8570 20516 8576 20528
rect 8242 20488 8576 20516
rect 8242 20485 8254 20488
rect 8196 20479 8254 20485
rect 8570 20476 8576 20488
rect 8628 20476 8634 20528
rect 9582 20476 9588 20528
rect 9640 20516 9646 20528
rect 9876 20516 9904 20547
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 13633 20587 13691 20593
rect 13633 20553 13645 20587
rect 13679 20584 13691 20587
rect 14734 20584 14740 20596
rect 13679 20556 14740 20584
rect 13679 20553 13691 20556
rect 13633 20547 13691 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 15378 20584 15384 20596
rect 15335 20556 15384 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 15654 20544 15660 20596
rect 15712 20544 15718 20596
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 15896 20556 17724 20584
rect 15896 20544 15902 20556
rect 9640 20488 9904 20516
rect 10220 20519 10278 20525
rect 9640 20476 9646 20488
rect 10220 20485 10232 20519
rect 10266 20516 10278 20519
rect 10318 20516 10324 20528
rect 10266 20488 10324 20516
rect 10266 20485 10278 20488
rect 10220 20479 10278 20485
rect 10318 20476 10324 20488
rect 10376 20476 10382 20528
rect 12520 20519 12578 20525
rect 12520 20485 12532 20519
rect 12566 20516 12578 20519
rect 12710 20516 12716 20528
rect 12566 20488 12716 20516
rect 12566 20485 12578 20488
rect 12520 20479 12578 20485
rect 12710 20476 12716 20488
rect 12768 20476 12774 20528
rect 15194 20516 15200 20528
rect 13924 20488 15200 20516
rect 7745 20451 7803 20457
rect 7745 20448 7757 20451
rect 7156 20420 7757 20448
rect 7156 20408 7162 20420
rect 7745 20417 7757 20420
rect 7791 20417 7803 20451
rect 7745 20411 7803 20417
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 9953 20451 10011 20457
rect 9953 20448 9965 20451
rect 9916 20420 9965 20448
rect 9916 20408 9922 20420
rect 9953 20417 9965 20420
rect 9999 20448 10011 20451
rect 11238 20448 11244 20460
rect 9999 20420 11244 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 11330 20408 11336 20460
rect 11388 20448 11394 20460
rect 13924 20457 13952 20488
rect 15194 20476 15200 20488
rect 15252 20516 15258 20528
rect 16206 20516 16212 20528
rect 15252 20488 16212 20516
rect 15252 20476 15258 20488
rect 16206 20476 16212 20488
rect 16264 20516 16270 20528
rect 16482 20516 16488 20528
rect 16264 20488 16488 20516
rect 16264 20476 16270 20488
rect 16482 20476 16488 20488
rect 16540 20516 16546 20528
rect 17589 20519 17647 20525
rect 17589 20516 17601 20519
rect 16540 20488 17601 20516
rect 16540 20476 16546 20488
rect 17589 20485 17601 20488
rect 17635 20485 17647 20519
rect 17589 20479 17647 20485
rect 12069 20451 12127 20457
rect 12069 20448 12081 20451
rect 11388 20420 12081 20448
rect 11388 20408 11394 20420
rect 12069 20417 12081 20420
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 13998 20408 14004 20460
rect 14056 20448 14062 20460
rect 14165 20451 14223 20457
rect 14165 20448 14177 20451
rect 14056 20420 14177 20448
rect 14056 20408 14062 20420
rect 14165 20417 14177 20420
rect 14211 20417 14223 20451
rect 14165 20411 14223 20417
rect 14458 20408 14464 20460
rect 14516 20448 14522 20460
rect 14734 20448 14740 20460
rect 14516 20420 14740 20448
rect 14516 20408 14522 20420
rect 14734 20408 14740 20420
rect 14792 20448 14798 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 14792 20420 15761 20448
rect 14792 20408 14798 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 3237 20383 3295 20389
rect 3237 20349 3249 20383
rect 3283 20349 3295 20383
rect 3237 20343 3295 20349
rect 4801 20383 4859 20389
rect 4801 20349 4813 20383
rect 4847 20349 4859 20383
rect 4801 20343 4859 20349
rect 3252 20244 3280 20343
rect 4816 20312 4844 20343
rect 6454 20340 6460 20392
rect 6512 20340 6518 20392
rect 6641 20383 6699 20389
rect 6641 20349 6653 20383
rect 6687 20380 6699 20383
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 6687 20352 7205 20380
rect 6687 20349 6699 20352
rect 6641 20343 6699 20349
rect 7193 20349 7205 20352
rect 7239 20349 7251 20383
rect 11256 20380 11284 20408
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 11256 20352 12265 20380
rect 7193 20343 7251 20349
rect 12253 20349 12265 20352
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 15562 20340 15568 20392
rect 15620 20380 15626 20392
rect 16022 20380 16028 20392
rect 15620 20352 16028 20380
rect 15620 20340 15626 20352
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 16316 20380 16344 20411
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16816 20420 16865 20448
rect 16816 20408 16822 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17218 20380 17224 20392
rect 16316 20352 17224 20380
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 17696 20380 17724 20556
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 20036 20556 20085 20584
rect 20036 20544 20042 20556
rect 20073 20553 20085 20556
rect 20119 20553 20131 20587
rect 20346 20584 20352 20596
rect 20073 20547 20131 20553
rect 20180 20556 20352 20584
rect 18966 20457 18972 20460
rect 18944 20451 18972 20457
rect 18944 20417 18956 20451
rect 18944 20411 18972 20417
rect 18966 20408 18972 20411
rect 19024 20408 19030 20460
rect 19794 20408 19800 20460
rect 19852 20408 19858 20460
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20180 20448 20208 20556
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 20533 20587 20591 20593
rect 20533 20553 20545 20587
rect 20579 20584 20591 20587
rect 21266 20584 21272 20596
rect 20579 20556 21272 20584
rect 20579 20553 20591 20556
rect 20533 20547 20591 20553
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 20714 20516 20720 20528
rect 20272 20488 20720 20516
rect 20272 20457 20300 20488
rect 20714 20476 20720 20488
rect 20772 20476 20778 20528
rect 20027 20420 20208 20448
rect 20257 20451 20315 20457
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20257 20417 20269 20451
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 18785 20383 18843 20389
rect 18785 20380 18797 20383
rect 17696 20352 18797 20380
rect 18785 20349 18797 20352
rect 18831 20349 18843 20383
rect 18785 20343 18843 20349
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20380 19119 20383
rect 19242 20380 19248 20392
rect 19107 20352 19248 20380
rect 19107 20349 19119 20352
rect 19061 20343 19119 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 19334 20340 19340 20392
rect 19392 20340 19398 20392
rect 4172 20284 4844 20312
rect 16485 20315 16543 20321
rect 4172 20256 4200 20284
rect 16485 20281 16497 20315
rect 16531 20312 16543 20315
rect 16942 20312 16948 20324
rect 16531 20284 16948 20312
rect 16531 20281 16543 20284
rect 16485 20275 16543 20281
rect 16942 20272 16948 20284
rect 17000 20272 17006 20324
rect 4154 20244 4160 20256
rect 3252 20216 4160 20244
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 11514 20204 11520 20256
rect 11572 20204 11578 20256
rect 15930 20204 15936 20256
rect 15988 20244 15994 20256
rect 16117 20247 16175 20253
rect 16117 20244 16129 20247
rect 15988 20216 16129 20244
rect 15988 20204 15994 20216
rect 16117 20213 16129 20216
rect 16163 20213 16175 20247
rect 16117 20207 16175 20213
rect 18141 20247 18199 20253
rect 18141 20213 18153 20247
rect 18187 20244 18199 20247
rect 20364 20244 20392 20411
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23658 20408 23664 20460
rect 23716 20408 23722 20460
rect 18187 20216 20392 20244
rect 18187 20213 18199 20216
rect 18141 20207 18199 20213
rect 22186 20204 22192 20256
rect 22244 20244 22250 20256
rect 23109 20247 23167 20253
rect 23109 20244 23121 20247
rect 22244 20216 23121 20244
rect 22244 20204 22250 20216
rect 23109 20213 23121 20216
rect 23155 20213 23167 20247
rect 23109 20207 23167 20213
rect 23474 20204 23480 20256
rect 23532 20204 23538 20256
rect 1104 20154 24012 20176
rect 1104 20102 1350 20154
rect 1402 20102 1414 20154
rect 1466 20102 1478 20154
rect 1530 20102 1542 20154
rect 1594 20102 1606 20154
rect 1658 20102 4350 20154
rect 4402 20102 4414 20154
rect 4466 20102 4478 20154
rect 4530 20102 4542 20154
rect 4594 20102 4606 20154
rect 4658 20102 7350 20154
rect 7402 20102 7414 20154
rect 7466 20102 7478 20154
rect 7530 20102 7542 20154
rect 7594 20102 7606 20154
rect 7658 20102 10350 20154
rect 10402 20102 10414 20154
rect 10466 20102 10478 20154
rect 10530 20102 10542 20154
rect 10594 20102 10606 20154
rect 10658 20102 13350 20154
rect 13402 20102 13414 20154
rect 13466 20102 13478 20154
rect 13530 20102 13542 20154
rect 13594 20102 13606 20154
rect 13658 20102 16350 20154
rect 16402 20102 16414 20154
rect 16466 20102 16478 20154
rect 16530 20102 16542 20154
rect 16594 20102 16606 20154
rect 16658 20102 19350 20154
rect 19402 20102 19414 20154
rect 19466 20102 19478 20154
rect 19530 20102 19542 20154
rect 19594 20102 19606 20154
rect 19658 20102 22350 20154
rect 22402 20102 22414 20154
rect 22466 20102 22478 20154
rect 22530 20102 22542 20154
rect 22594 20102 22606 20154
rect 22658 20102 24012 20154
rect 1104 20080 24012 20102
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 7377 20043 7435 20049
rect 7377 20040 7389 20043
rect 7248 20012 7389 20040
rect 7248 20000 7254 20012
rect 7377 20009 7389 20012
rect 7423 20009 7435 20043
rect 7377 20003 7435 20009
rect 8754 20000 8760 20052
rect 8812 20040 8818 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8812 20012 8953 20040
rect 8812 20000 8818 20012
rect 8941 20009 8953 20012
rect 8987 20009 8999 20043
rect 8941 20003 8999 20009
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 10137 20043 10195 20049
rect 10137 20040 10149 20043
rect 9732 20012 10149 20040
rect 9732 20000 9738 20012
rect 10137 20009 10149 20012
rect 10183 20009 10195 20043
rect 10137 20003 10195 20009
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11756 20012 11897 20040
rect 11756 20000 11762 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 13964 20012 14381 20040
rect 13964 20000 13970 20012
rect 14369 20009 14381 20012
rect 14415 20009 14427 20043
rect 14369 20003 14427 20009
rect 16114 20000 16120 20052
rect 16172 20000 16178 20052
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19242 20040 19248 20052
rect 18932 20012 19248 20040
rect 18932 20000 18938 20012
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 19429 20043 19487 20049
rect 19429 20009 19441 20043
rect 19475 20040 19487 20043
rect 19702 20040 19708 20052
rect 19475 20012 19708 20040
rect 19475 20009 19487 20012
rect 19429 20003 19487 20009
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 11514 19972 11520 19984
rect 10612 19944 11520 19972
rect 9490 19864 9496 19916
rect 9548 19864 9554 19916
rect 10612 19913 10640 19944
rect 11514 19932 11520 19944
rect 11572 19932 11578 19984
rect 10597 19907 10655 19913
rect 10597 19873 10609 19907
rect 10643 19873 10655 19907
rect 10597 19867 10655 19873
rect 10778 19864 10784 19916
rect 10836 19864 10842 19916
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 11204 19876 12112 19904
rect 11204 19864 11210 19876
rect 6638 19796 6644 19848
rect 6696 19836 6702 19848
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 6696 19808 7205 19836
rect 6696 19796 6702 19808
rect 7193 19805 7205 19808
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 9398 19836 9404 19848
rect 9355 19808 9404 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 9398 19796 9404 19808
rect 9456 19836 9462 19848
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 9456 19808 10517 19836
rect 9456 19796 9462 19808
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 12084 19845 12112 19876
rect 14366 19864 14372 19916
rect 14424 19904 14430 19916
rect 14921 19907 14979 19913
rect 14921 19904 14933 19907
rect 14424 19876 14933 19904
rect 14424 19864 14430 19876
rect 14921 19873 14933 19876
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15436 19876 15761 19904
rect 15436 19864 15442 19876
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 15749 19867 15807 19873
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 17678 19904 17684 19916
rect 17552 19876 17684 19904
rect 17552 19864 17558 19876
rect 17678 19864 17684 19876
rect 17736 19904 17742 19916
rect 17773 19907 17831 19913
rect 17773 19904 17785 19907
rect 17736 19876 17785 19904
rect 17736 19864 17742 19876
rect 17773 19873 17785 19876
rect 17819 19873 17831 19907
rect 17773 19867 17831 19873
rect 18693 19907 18751 19913
rect 18693 19873 18705 19907
rect 18739 19904 18751 19907
rect 18966 19904 18972 19916
rect 18739 19876 18972 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 11609 19839 11667 19845
rect 11609 19836 11621 19839
rect 11296 19808 11621 19836
rect 11296 19796 11302 19808
rect 11609 19805 11621 19808
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 14734 19796 14740 19848
rect 14792 19796 14798 19848
rect 15930 19796 15936 19848
rect 15988 19796 15994 19848
rect 16206 19796 16212 19848
rect 16264 19836 16270 19848
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 16264 19808 17049 19836
rect 16264 19796 16270 19808
rect 17037 19805 17049 19808
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19836 17647 19839
rect 18598 19836 18604 19848
rect 17635 19808 18604 19836
rect 17635 19805 17647 19808
rect 17589 19799 17647 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19208 19808 19257 19836
rect 19208 19796 19214 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 22830 19796 22836 19848
rect 22888 19796 22894 19848
rect 22925 19839 22983 19845
rect 22925 19805 22937 19839
rect 22971 19805 22983 19839
rect 22925 19799 22983 19805
rect 22738 19728 22744 19780
rect 22796 19768 22802 19780
rect 22940 19768 22968 19799
rect 23014 19796 23020 19848
rect 23072 19836 23078 19848
rect 23385 19839 23443 19845
rect 23385 19836 23397 19839
rect 23072 19808 23397 19836
rect 23072 19796 23078 19808
rect 23385 19805 23397 19808
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 23750 19836 23756 19848
rect 23707 19808 23756 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 22796 19740 22968 19768
rect 22796 19728 22802 19740
rect 9398 19660 9404 19712
rect 9456 19660 9462 19712
rect 14829 19703 14887 19709
rect 14829 19669 14841 19703
rect 14875 19700 14887 19703
rect 15197 19703 15255 19709
rect 15197 19700 15209 19703
rect 14875 19672 15209 19700
rect 14875 19669 14887 19672
rect 14829 19663 14887 19669
rect 15197 19669 15209 19672
rect 15243 19669 15255 19703
rect 15197 19663 15255 19669
rect 17681 19703 17739 19709
rect 17681 19669 17693 19703
rect 17727 19700 17739 19703
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 17727 19672 18061 19700
rect 17727 19669 17739 19672
rect 17681 19663 17739 19669
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18049 19663 18107 19669
rect 21818 19660 21824 19712
rect 21876 19700 21882 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 21876 19672 22661 19700
rect 21876 19660 21882 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 22649 19663 22707 19669
rect 23106 19660 23112 19712
rect 23164 19660 23170 19712
rect 23198 19660 23204 19712
rect 23256 19660 23262 19712
rect 23477 19703 23535 19709
rect 23477 19669 23489 19703
rect 23523 19700 23535 19703
rect 23658 19700 23664 19712
rect 23523 19672 23664 19700
rect 23523 19669 23535 19672
rect 23477 19663 23535 19669
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 1104 19610 24164 19632
rect 1104 19558 2850 19610
rect 2902 19558 2914 19610
rect 2966 19558 2978 19610
rect 3030 19558 3042 19610
rect 3094 19558 3106 19610
rect 3158 19558 5850 19610
rect 5902 19558 5914 19610
rect 5966 19558 5978 19610
rect 6030 19558 6042 19610
rect 6094 19558 6106 19610
rect 6158 19558 8850 19610
rect 8902 19558 8914 19610
rect 8966 19558 8978 19610
rect 9030 19558 9042 19610
rect 9094 19558 9106 19610
rect 9158 19558 11850 19610
rect 11902 19558 11914 19610
rect 11966 19558 11978 19610
rect 12030 19558 12042 19610
rect 12094 19558 12106 19610
rect 12158 19558 14850 19610
rect 14902 19558 14914 19610
rect 14966 19558 14978 19610
rect 15030 19558 15042 19610
rect 15094 19558 15106 19610
rect 15158 19558 17850 19610
rect 17902 19558 17914 19610
rect 17966 19558 17978 19610
rect 18030 19558 18042 19610
rect 18094 19558 18106 19610
rect 18158 19558 20850 19610
rect 20902 19558 20914 19610
rect 20966 19558 20978 19610
rect 21030 19558 21042 19610
rect 21094 19558 21106 19610
rect 21158 19558 23850 19610
rect 23902 19558 23914 19610
rect 23966 19558 23978 19610
rect 24030 19558 24042 19610
rect 24094 19558 24106 19610
rect 24158 19558 24164 19610
rect 1104 19536 24164 19558
rect 7929 19499 7987 19505
rect 7929 19496 7941 19499
rect 1688 19468 7941 19496
rect 1688 19369 1716 19468
rect 7929 19465 7941 19468
rect 7975 19465 7987 19499
rect 7929 19459 7987 19465
rect 9398 19456 9404 19508
rect 9456 19456 9462 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11606 19496 11612 19508
rect 11563 19468 11612 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 13320 19468 13461 19496
rect 13320 19456 13326 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 13449 19459 13507 19465
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15286 19496 15292 19508
rect 15243 19468 15292 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 16942 19496 16948 19508
rect 16715 19468 16948 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 5626 19388 5632 19440
rect 5684 19428 5690 19440
rect 5684 19400 8156 19428
rect 5684 19388 5690 19400
rect 3510 19369 3516 19372
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 3504 19323 3516 19369
rect 3510 19320 3516 19323
rect 3568 19320 3574 19372
rect 4632 19332 6040 19360
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19261 3295 19295
rect 3237 19255 3295 19261
rect 1210 19116 1216 19168
rect 1268 19156 1274 19168
rect 1489 19159 1547 19165
rect 1489 19156 1501 19159
rect 1268 19128 1501 19156
rect 1268 19116 1274 19128
rect 1489 19125 1501 19128
rect 1535 19125 1547 19159
rect 3252 19156 3280 19255
rect 4632 19233 4660 19332
rect 5258 19252 5264 19304
rect 5316 19252 5322 19304
rect 6012 19301 6040 19332
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 6696 19332 6745 19360
rect 6696 19320 6702 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 6825 19363 6883 19369
rect 6825 19329 6837 19363
rect 6871 19360 6883 19363
rect 7006 19360 7012 19372
rect 6871 19332 7012 19360
rect 6871 19329 6883 19332
rect 6825 19323 6883 19329
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 8128 19369 8156 19400
rect 23106 19388 23112 19440
rect 23164 19388 23170 19440
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 9674 19320 9680 19372
rect 9732 19360 9738 19372
rect 10597 19363 10655 19369
rect 10597 19360 10609 19363
rect 9732 19332 10609 19360
rect 9732 19320 9738 19332
rect 10597 19329 10609 19332
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11112 19332 11713 19360
rect 11112 19320 11118 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 13357 19363 13415 19369
rect 13357 19329 13369 19363
rect 13403 19360 13415 19363
rect 13817 19363 13875 19369
rect 13817 19360 13829 19363
rect 13403 19332 13829 19360
rect 13403 19329 13415 19332
rect 13357 19323 13415 19329
rect 13817 19329 13829 19332
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 13906 19320 13912 19372
rect 13964 19360 13970 19372
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 13964 19332 15393 19360
rect 13964 19320 13970 19332
rect 15381 19329 15393 19332
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 16264 19332 16313 19360
rect 16264 19320 16270 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 17678 19360 17684 19372
rect 16899 19332 17684 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 17770 19320 17776 19372
rect 17828 19320 17834 19372
rect 20714 19320 20720 19372
rect 20772 19320 20778 19372
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21324 19332 21833 19360
rect 21324 19320 21330 19332
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 23124 19360 23152 19388
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 23124 19332 23397 19360
rect 21821 19323 21879 19329
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 5997 19295 6055 19301
rect 5997 19261 6009 19295
rect 6043 19292 6055 19295
rect 6086 19292 6092 19304
rect 6043 19264 6092 19292
rect 6043 19261 6055 19264
rect 5997 19255 6055 19261
rect 6086 19252 6092 19264
rect 6144 19252 6150 19304
rect 6546 19252 6552 19304
rect 6604 19292 6610 19304
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6604 19264 6929 19292
rect 6604 19252 6610 19264
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 6917 19255 6975 19261
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7745 19295 7803 19301
rect 7745 19292 7757 19295
rect 7156 19264 7757 19292
rect 7156 19252 7162 19264
rect 7745 19261 7757 19264
rect 7791 19261 7803 19295
rect 7745 19255 7803 19261
rect 9306 19252 9312 19304
rect 9364 19292 9370 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9364 19264 9965 19292
rect 9364 19252 9370 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 10686 19252 10692 19304
rect 10744 19252 10750 19304
rect 10870 19252 10876 19304
rect 10928 19292 10934 19304
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 10928 19264 11253 19292
rect 10928 19252 10934 19264
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 11241 19255 11299 19261
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 4617 19227 4675 19233
rect 4617 19193 4629 19227
rect 4663 19193 4675 19227
rect 4617 19187 4675 19193
rect 6454 19184 6460 19236
rect 6512 19224 6518 19236
rect 10226 19224 10232 19236
rect 6512 19196 10232 19224
rect 6512 19184 6518 19196
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 10704 19224 10732 19252
rect 12342 19224 12348 19236
rect 10704 19196 12348 19224
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 13648 19224 13676 19255
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14240 19264 14381 19292
rect 14240 19252 14246 19264
rect 14369 19261 14381 19264
rect 14415 19261 14427 19295
rect 14369 19255 14427 19261
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19292 18475 19295
rect 18782 19292 18788 19304
rect 18463 19264 18788 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19292 19671 19295
rect 19794 19292 19800 19304
rect 19659 19264 19800 19292
rect 19659 19261 19671 19264
rect 19613 19255 19671 19261
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 22465 19295 22523 19301
rect 22465 19261 22477 19295
rect 22511 19292 22523 19295
rect 22922 19292 22928 19304
rect 22511 19264 22928 19292
rect 22511 19261 22523 19264
rect 22465 19255 22523 19261
rect 22922 19252 22928 19264
rect 22980 19252 22986 19304
rect 23106 19252 23112 19304
rect 23164 19252 23170 19304
rect 13722 19224 13728 19236
rect 13648 19196 13728 19224
rect 13722 19184 13728 19196
rect 13780 19224 13786 19236
rect 15654 19224 15660 19236
rect 13780 19196 15660 19224
rect 13780 19184 13786 19196
rect 15654 19184 15660 19196
rect 15712 19184 15718 19236
rect 19886 19184 19892 19236
rect 19944 19224 19950 19236
rect 23474 19224 23480 19236
rect 19944 19196 23480 19224
rect 19944 19184 19950 19196
rect 23474 19184 23480 19196
rect 23532 19184 23538 19236
rect 4154 19156 4160 19168
rect 3252 19128 4160 19156
rect 1489 19119 1547 19125
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4706 19116 4712 19168
rect 4764 19116 4770 19168
rect 5442 19116 5448 19168
rect 5500 19116 5506 19168
rect 6362 19116 6368 19168
rect 6420 19116 6426 19168
rect 7190 19116 7196 19168
rect 7248 19116 7254 19168
rect 10686 19116 10692 19168
rect 10744 19116 10750 19168
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 12989 19159 13047 19165
rect 12989 19156 13001 19159
rect 12768 19128 13001 19156
rect 12768 19116 12774 19128
rect 12989 19125 13001 19128
rect 13035 19125 13047 19159
rect 12989 19119 13047 19125
rect 16114 19116 16120 19168
rect 16172 19116 16178 19168
rect 19702 19116 19708 19168
rect 19760 19156 19766 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19760 19128 20177 19156
rect 19760 19116 19766 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20165 19119 20223 19125
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 20496 19128 20545 19156
rect 20496 19116 20502 19128
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 20533 19119 20591 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22557 19159 22615 19165
rect 22557 19156 22569 19159
rect 22152 19128 22569 19156
rect 22152 19116 22158 19128
rect 22557 19125 22569 19128
rect 22603 19125 22615 19159
rect 22557 19119 22615 19125
rect 23566 19116 23572 19168
rect 23624 19116 23630 19168
rect 1104 19066 24012 19088
rect 1104 19014 1350 19066
rect 1402 19014 1414 19066
rect 1466 19014 1478 19066
rect 1530 19014 1542 19066
rect 1594 19014 1606 19066
rect 1658 19014 4350 19066
rect 4402 19014 4414 19066
rect 4466 19014 4478 19066
rect 4530 19014 4542 19066
rect 4594 19014 4606 19066
rect 4658 19014 7350 19066
rect 7402 19014 7414 19066
rect 7466 19014 7478 19066
rect 7530 19014 7542 19066
rect 7594 19014 7606 19066
rect 7658 19014 10350 19066
rect 10402 19014 10414 19066
rect 10466 19014 10478 19066
rect 10530 19014 10542 19066
rect 10594 19014 10606 19066
rect 10658 19014 13350 19066
rect 13402 19014 13414 19066
rect 13466 19014 13478 19066
rect 13530 19014 13542 19066
rect 13594 19014 13606 19066
rect 13658 19014 16350 19066
rect 16402 19014 16414 19066
rect 16466 19014 16478 19066
rect 16530 19014 16542 19066
rect 16594 19014 16606 19066
rect 16658 19014 19350 19066
rect 19402 19014 19414 19066
rect 19466 19014 19478 19066
rect 19530 19014 19542 19066
rect 19594 19014 19606 19066
rect 19658 19014 22350 19066
rect 22402 19014 22414 19066
rect 22466 19014 22478 19066
rect 22530 19014 22542 19066
rect 22594 19014 22606 19066
rect 22658 19014 24012 19066
rect 1104 18992 24012 19014
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 3510 18952 3516 18964
rect 3467 18924 3516 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 5169 18955 5227 18961
rect 5169 18921 5181 18955
rect 5215 18952 5227 18955
rect 5626 18952 5632 18964
rect 5215 18924 5632 18952
rect 5215 18921 5227 18924
rect 5169 18915 5227 18921
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 7098 18912 7104 18964
rect 7156 18912 7162 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 21358 18952 21364 18964
rect 16172 18924 21364 18952
rect 16172 18912 16178 18924
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 1627 18856 2774 18884
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 2746 18816 2774 18856
rect 4801 18819 4859 18825
rect 2746 18788 4568 18816
rect 382 18708 388 18760
rect 440 18748 446 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 440 18720 1409 18748
rect 440 18708 446 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 3602 18708 3608 18760
rect 3660 18708 3666 18760
rect 4540 18757 4568 18788
rect 4801 18785 4813 18819
rect 4847 18816 4859 18819
rect 4847 18788 5212 18816
rect 4847 18785 4859 18788
rect 4801 18779 4859 18785
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18748 4031 18751
rect 4525 18751 4583 18757
rect 4019 18720 4200 18748
rect 4019 18717 4031 18720
rect 3973 18711 4031 18717
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 4172 18621 4200 18720
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 5074 18748 5080 18760
rect 4571 18720 5080 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 4706 18680 4712 18692
rect 4663 18652 4712 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 4706 18640 4712 18652
rect 4764 18640 4770 18692
rect 4157 18615 4215 18621
rect 4157 18581 4169 18615
rect 4203 18581 4215 18615
rect 5184 18612 5212 18788
rect 5258 18776 5264 18828
rect 5316 18816 5322 18828
rect 5951 18819 6009 18825
rect 5951 18816 5963 18819
rect 5316 18788 5963 18816
rect 5316 18776 5322 18788
rect 5951 18785 5963 18788
rect 5997 18785 6009 18819
rect 5951 18779 6009 18785
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 6270 18776 6276 18828
rect 6328 18816 6334 18828
rect 6365 18819 6423 18825
rect 6365 18816 6377 18819
rect 6328 18788 6377 18816
rect 6328 18776 6334 18788
rect 6365 18785 6377 18788
rect 6411 18816 6423 18819
rect 6730 18816 6736 18828
rect 6411 18788 6736 18816
rect 6411 18785 6423 18788
rect 6365 18779 6423 18785
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 6825 18819 6883 18825
rect 6825 18785 6837 18819
rect 6871 18816 6883 18819
rect 7116 18816 7144 18912
rect 12989 18887 13047 18893
rect 12989 18853 13001 18887
rect 13035 18853 13047 18887
rect 12989 18847 13047 18853
rect 19245 18887 19303 18893
rect 19245 18853 19257 18887
rect 19291 18853 19303 18887
rect 19245 18847 19303 18853
rect 6871 18788 7144 18816
rect 8481 18819 8539 18825
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 9674 18816 9680 18828
rect 8527 18788 9680 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10226 18776 10232 18828
rect 10284 18816 10290 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 10284 18788 10425 18816
rect 10284 18776 10290 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 10413 18779 10471 18785
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7009 18751 7067 18757
rect 7009 18748 7021 18751
rect 6972 18720 7021 18748
rect 6972 18708 6978 18720
rect 7009 18717 7021 18720
rect 7055 18717 7067 18751
rect 9490 18748 9496 18760
rect 7009 18711 7067 18717
rect 7116 18720 9496 18748
rect 7116 18612 7144 18720
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 9582 18708 9588 18760
rect 9640 18708 9646 18760
rect 9692 18748 9720 18776
rect 11517 18751 11575 18757
rect 11517 18748 11529 18751
rect 9692 18720 11529 18748
rect 11517 18717 11529 18720
rect 11563 18748 11575 18751
rect 11698 18748 11704 18760
rect 11563 18720 11704 18748
rect 11563 18717 11575 18720
rect 11517 18711 11575 18717
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 12713 18751 12771 18757
rect 12713 18717 12725 18751
rect 12759 18748 12771 18751
rect 13004 18748 13032 18847
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 13814 18816 13820 18828
rect 13679 18788 13820 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 15344 18788 15669 18816
rect 15344 18776 15350 18788
rect 15657 18785 15669 18788
rect 15703 18785 15715 18819
rect 15657 18779 15715 18785
rect 12759 18720 13032 18748
rect 12759 18717 12771 18720
rect 12713 18711 12771 18717
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 13320 18720 13369 18748
rect 13320 18708 13326 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 7742 18640 7748 18692
rect 7800 18680 7806 18692
rect 8214 18683 8272 18689
rect 8214 18680 8226 18683
rect 7800 18652 8226 18680
rect 7800 18640 7806 18652
rect 8214 18649 8226 18652
rect 8260 18649 8272 18683
rect 8214 18643 8272 18649
rect 8662 18640 8668 18692
rect 8720 18680 8726 18692
rect 10229 18683 10287 18689
rect 10229 18680 10241 18683
rect 8720 18652 10241 18680
rect 8720 18640 8726 18652
rect 10229 18649 10241 18652
rect 10275 18649 10287 18683
rect 10229 18643 10287 18649
rect 10321 18683 10379 18689
rect 10321 18649 10333 18683
rect 10367 18680 10379 18683
rect 10686 18680 10692 18692
rect 10367 18652 10692 18680
rect 10367 18649 10379 18652
rect 10321 18643 10379 18649
rect 10686 18640 10692 18652
rect 10744 18640 10750 18692
rect 10781 18683 10839 18689
rect 10781 18649 10793 18683
rect 10827 18680 10839 18683
rect 10962 18680 10968 18692
rect 10827 18652 10968 18680
rect 10827 18649 10839 18652
rect 10781 18643 10839 18649
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 13372 18680 13400 18711
rect 14458 18708 14464 18760
rect 14516 18748 14522 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14516 18720 14657 18748
rect 14516 18708 14522 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 15013 18751 15071 18757
rect 15013 18717 15025 18751
rect 15059 18748 15071 18751
rect 15378 18748 15384 18760
rect 15059 18720 15384 18748
rect 15059 18717 15071 18720
rect 15013 18711 15071 18717
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18748 15531 18751
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15519 18720 16405 18748
rect 15519 18717 15531 18720
rect 15473 18711 15531 18717
rect 16393 18717 16405 18720
rect 16439 18748 16451 18751
rect 17402 18748 17408 18760
rect 16439 18720 17408 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 18598 18708 18604 18760
rect 18656 18708 18662 18760
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 19260 18748 19288 18847
rect 19702 18776 19708 18828
rect 19760 18776 19766 18828
rect 19812 18825 19840 18924
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 22557 18955 22615 18961
rect 22557 18921 22569 18955
rect 22603 18952 22615 18955
rect 22830 18952 22836 18964
rect 22603 18924 22836 18952
rect 22603 18921 22615 18924
rect 22557 18915 22615 18921
rect 22830 18912 22836 18924
rect 22888 18912 22894 18964
rect 21545 18887 21603 18893
rect 21545 18853 21557 18887
rect 21591 18884 21603 18887
rect 22922 18884 22928 18896
rect 21591 18856 22928 18884
rect 21591 18853 21603 18856
rect 21545 18847 21603 18853
rect 22922 18844 22928 18856
rect 22980 18844 22986 18896
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 20162 18776 20168 18828
rect 20220 18776 20226 18828
rect 22005 18819 22063 18825
rect 22005 18785 22017 18819
rect 22051 18785 22063 18819
rect 22005 18779 22063 18785
rect 18739 18720 19288 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19392 18720 19625 18748
rect 19392 18708 19398 18720
rect 19613 18717 19625 18720
rect 19659 18748 19671 18751
rect 19886 18748 19892 18760
rect 19659 18720 19892 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 20438 18757 20444 18760
rect 20432 18748 20444 18757
rect 20399 18720 20444 18748
rect 20432 18711 20444 18720
rect 20438 18708 20444 18711
rect 20496 18708 20502 18760
rect 22020 18748 22048 18779
rect 22094 18776 22100 18828
rect 22152 18776 22158 18828
rect 22370 18816 22376 18828
rect 22204 18788 22376 18816
rect 22204 18748 22232 18788
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 22020 18720 22232 18748
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23201 18751 23259 18757
rect 23201 18748 23213 18751
rect 22796 18720 23213 18748
rect 22796 18708 22802 18720
rect 23201 18717 23213 18720
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18717 23443 18751
rect 23385 18711 23443 18717
rect 16660 18683 16718 18689
rect 13372 18652 14688 18680
rect 14660 18624 14688 18652
rect 16660 18649 16672 18683
rect 16706 18680 16718 18683
rect 16850 18680 16856 18692
rect 16706 18652 16856 18680
rect 16706 18649 16718 18652
rect 16660 18643 16718 18649
rect 16850 18640 16856 18652
rect 16908 18640 16914 18692
rect 18782 18680 18788 18692
rect 17788 18652 18788 18680
rect 5184 18584 7144 18612
rect 4157 18575 4215 18581
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 8941 18615 8999 18621
rect 8941 18612 8953 18615
rect 8812 18584 8953 18612
rect 8812 18572 8818 18584
rect 8941 18581 8953 18584
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 9861 18615 9919 18621
rect 9861 18612 9873 18615
rect 9364 18584 9873 18612
rect 9364 18572 9370 18584
rect 9861 18581 9873 18584
rect 9907 18581 9919 18615
rect 9861 18575 9919 18581
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 13449 18615 13507 18621
rect 13449 18581 13461 18615
rect 13495 18612 13507 18615
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13495 18584 14105 18612
rect 13495 18581 13507 18584
rect 13449 18575 13507 18581
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 14642 18572 14648 18624
rect 14700 18572 14706 18624
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 14829 18615 14887 18621
rect 14829 18612 14841 18615
rect 14792 18584 14841 18612
rect 14792 18572 14798 18584
rect 14829 18581 14841 18584
rect 14875 18581 14887 18615
rect 14829 18575 14887 18581
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 17788 18621 17816 18652
rect 18782 18640 18788 18652
rect 18840 18640 18846 18692
rect 19978 18640 19984 18692
rect 20036 18680 20042 18692
rect 23400 18680 23428 18711
rect 20036 18652 23428 18680
rect 20036 18640 20042 18652
rect 16301 18615 16359 18621
rect 16301 18612 16313 18615
rect 16080 18584 16313 18612
rect 16080 18572 16086 18584
rect 16301 18581 16313 18584
rect 16347 18581 16359 18615
rect 16301 18575 16359 18581
rect 17773 18615 17831 18621
rect 17773 18581 17785 18615
rect 17819 18581 17831 18615
rect 17773 18575 17831 18581
rect 17957 18615 18015 18621
rect 17957 18581 17969 18615
rect 18003 18612 18015 18615
rect 18230 18612 18236 18624
rect 18003 18584 18236 18612
rect 18003 18581 18015 18584
rect 17957 18575 18015 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 20254 18612 20260 18624
rect 18923 18584 20260 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22189 18615 22247 18621
rect 22189 18612 22201 18615
rect 22152 18584 22201 18612
rect 22152 18572 22158 18584
rect 22189 18581 22201 18584
rect 22235 18612 22247 18615
rect 22278 18612 22284 18624
rect 22235 18584 22284 18612
rect 22235 18581 22247 18584
rect 22189 18575 22247 18581
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22649 18615 22707 18621
rect 22649 18581 22661 18615
rect 22695 18612 22707 18615
rect 22738 18612 22744 18624
rect 22695 18584 22744 18612
rect 22695 18581 22707 18584
rect 22649 18575 22707 18581
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 23569 18615 23627 18621
rect 23569 18581 23581 18615
rect 23615 18612 23627 18615
rect 24302 18612 24308 18624
rect 23615 18584 24308 18612
rect 23615 18581 23627 18584
rect 23569 18575 23627 18581
rect 24302 18572 24308 18584
rect 24360 18572 24366 18624
rect 1104 18522 24164 18544
rect 1104 18470 2850 18522
rect 2902 18470 2914 18522
rect 2966 18470 2978 18522
rect 3030 18470 3042 18522
rect 3094 18470 3106 18522
rect 3158 18470 5850 18522
rect 5902 18470 5914 18522
rect 5966 18470 5978 18522
rect 6030 18470 6042 18522
rect 6094 18470 6106 18522
rect 6158 18470 8850 18522
rect 8902 18470 8914 18522
rect 8966 18470 8978 18522
rect 9030 18470 9042 18522
rect 9094 18470 9106 18522
rect 9158 18470 11850 18522
rect 11902 18470 11914 18522
rect 11966 18470 11978 18522
rect 12030 18470 12042 18522
rect 12094 18470 12106 18522
rect 12158 18470 14850 18522
rect 14902 18470 14914 18522
rect 14966 18470 14978 18522
rect 15030 18470 15042 18522
rect 15094 18470 15106 18522
rect 15158 18470 17850 18522
rect 17902 18470 17914 18522
rect 17966 18470 17978 18522
rect 18030 18470 18042 18522
rect 18094 18470 18106 18522
rect 18158 18470 20850 18522
rect 20902 18470 20914 18522
rect 20966 18470 20978 18522
rect 21030 18470 21042 18522
rect 21094 18470 21106 18522
rect 21158 18470 23850 18522
rect 23902 18470 23914 18522
rect 23966 18470 23978 18522
rect 24030 18470 24042 18522
rect 24094 18470 24106 18522
rect 24158 18470 24164 18522
rect 1104 18448 24164 18470
rect 3602 18368 3608 18420
rect 3660 18408 3666 18420
rect 4617 18411 4675 18417
rect 4617 18408 4629 18411
rect 3660 18380 4629 18408
rect 3660 18368 3666 18380
rect 4617 18377 4629 18380
rect 4663 18377 4675 18411
rect 4617 18371 4675 18377
rect 4985 18411 5043 18417
rect 4985 18377 4997 18411
rect 5031 18408 5043 18411
rect 5442 18408 5448 18420
rect 5031 18380 5448 18408
rect 5031 18377 5043 18380
rect 4985 18371 5043 18377
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 6733 18411 6791 18417
rect 6733 18377 6745 18411
rect 6779 18408 6791 18411
rect 7190 18408 7196 18420
rect 6779 18380 7196 18408
rect 6779 18377 6791 18380
rect 6733 18371 6791 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 8754 18368 8760 18420
rect 8812 18368 8818 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18377 9551 18411
rect 9493 18371 9551 18377
rect 3412 18343 3470 18349
rect 3412 18309 3424 18343
rect 3458 18340 3470 18343
rect 3786 18340 3792 18352
rect 3458 18312 3792 18340
rect 3458 18309 3470 18312
rect 3412 18303 3470 18309
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 5074 18300 5080 18352
rect 5132 18340 5138 18352
rect 6638 18340 6644 18352
rect 5132 18312 6644 18340
rect 5132 18300 5138 18312
rect 6638 18300 6644 18312
rect 6696 18340 6702 18352
rect 6825 18343 6883 18349
rect 6825 18340 6837 18343
rect 6696 18312 6837 18340
rect 6696 18300 6702 18312
rect 6825 18309 6837 18312
rect 6871 18309 6883 18343
rect 6825 18303 6883 18309
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 7285 18343 7343 18349
rect 7285 18340 7297 18343
rect 7064 18312 7297 18340
rect 7064 18300 7070 18312
rect 7285 18309 7297 18312
rect 7331 18309 7343 18343
rect 7285 18303 7343 18309
rect 8662 18300 8668 18352
rect 8720 18340 8726 18352
rect 8849 18343 8907 18349
rect 8849 18340 8861 18343
rect 8720 18312 8861 18340
rect 8720 18300 8726 18312
rect 8849 18309 8861 18312
rect 8895 18309 8907 18343
rect 9508 18340 9536 18371
rect 10870 18368 10876 18420
rect 10928 18408 10934 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10928 18380 10977 18408
rect 10928 18368 10934 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 11149 18411 11207 18417
rect 11149 18377 11161 18411
rect 11195 18377 11207 18411
rect 11149 18371 11207 18377
rect 13449 18411 13507 18417
rect 13449 18377 13461 18411
rect 13495 18408 13507 18411
rect 14458 18408 14464 18420
rect 13495 18380 14464 18408
rect 13495 18377 13507 18380
rect 13449 18371 13507 18377
rect 9830 18343 9888 18349
rect 9830 18340 9842 18343
rect 9508 18312 9842 18340
rect 8849 18303 8907 18309
rect 9830 18309 9842 18312
rect 9876 18309 9888 18343
rect 9830 18303 9888 18309
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 11164 18340 11192 18371
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 14700 18380 15332 18408
rect 14700 18368 14706 18380
rect 10284 18312 11192 18340
rect 12336 18343 12394 18349
rect 10284 18300 10290 18312
rect 12336 18309 12348 18343
rect 12382 18340 12394 18343
rect 12526 18340 12532 18352
rect 12382 18312 12532 18340
rect 12382 18309 12394 18312
rect 12336 18303 12394 18309
rect 12526 18300 12532 18312
rect 12584 18300 12590 18352
rect 15304 18340 15332 18380
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 15565 18411 15623 18417
rect 15565 18408 15577 18411
rect 15436 18380 15577 18408
rect 15436 18368 15442 18380
rect 15565 18377 15577 18380
rect 15611 18377 15623 18411
rect 15565 18371 15623 18377
rect 16022 18368 16028 18420
rect 16080 18368 16086 18420
rect 18506 18368 18512 18420
rect 18564 18408 18570 18420
rect 18564 18380 19932 18408
rect 18564 18368 18570 18380
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 15304 18312 15945 18340
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 19702 18340 19708 18352
rect 15933 18303 15991 18309
rect 19536 18312 19708 18340
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6362 18272 6368 18284
rect 5859 18244 6368 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 6512 18244 6592 18272
rect 6512 18232 6518 18244
rect 3145 18207 3203 18213
rect 3145 18173 3157 18207
rect 3191 18173 3203 18207
rect 3145 18167 3203 18173
rect 3160 18068 3188 18167
rect 5166 18164 5172 18216
rect 5224 18204 5230 18216
rect 6564 18213 6592 18244
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 9306 18232 9312 18284
rect 9364 18232 9370 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9674 18272 9680 18284
rect 9631 18244 9680 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 11146 18232 11152 18284
rect 11204 18272 11210 18284
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 11204 18244 11345 18272
rect 11204 18232 11210 18244
rect 11333 18241 11345 18244
rect 11379 18241 11391 18275
rect 11333 18235 11391 18241
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 12710 18272 12716 18284
rect 11839 18244 12716 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 14458 18281 14464 18284
rect 14436 18275 14464 18281
rect 14436 18241 14448 18275
rect 14436 18235 14464 18241
rect 14458 18232 14464 18235
rect 14516 18232 14522 18284
rect 14550 18232 14556 18284
rect 14608 18232 14614 18284
rect 15838 18272 15844 18284
rect 15120 18244 15844 18272
rect 6549 18207 6607 18213
rect 5224 18176 6500 18204
rect 5224 18164 5230 18176
rect 4525 18139 4583 18145
rect 4525 18105 4537 18139
rect 4571 18136 4583 18139
rect 5258 18136 5264 18148
rect 4571 18108 5264 18136
rect 4571 18105 4583 18108
rect 4525 18099 4583 18105
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 6472 18136 6500 18176
rect 6549 18173 6561 18207
rect 6595 18173 6607 18207
rect 6549 18167 6607 18173
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 6972 18176 7849 18204
rect 6972 18164 6978 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 7837 18167 7895 18173
rect 8128 18176 8953 18204
rect 8128 18145 8156 18176
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 11756 18176 12081 18204
rect 11756 18164 11762 18176
rect 12069 18173 12081 18176
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 13633 18207 13691 18213
rect 13633 18173 13645 18207
rect 13679 18204 13691 18207
rect 13906 18204 13912 18216
rect 13679 18176 13912 18204
rect 13679 18173 13691 18176
rect 13633 18167 13691 18173
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 15120 18204 15148 18244
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 16666 18232 16672 18284
rect 16724 18232 16730 18284
rect 18782 18232 18788 18284
rect 18840 18232 18846 18284
rect 19536 18281 19564 18312
rect 19702 18300 19708 18312
rect 19760 18300 19766 18352
rect 19904 18340 19932 18380
rect 19978 18368 19984 18420
rect 20036 18368 20042 18420
rect 21453 18411 21511 18417
rect 21453 18377 21465 18411
rect 21499 18408 21511 18411
rect 22646 18408 22652 18420
rect 21499 18380 22652 18408
rect 21499 18377 21511 18380
rect 21453 18371 21511 18377
rect 22646 18368 22652 18380
rect 22704 18368 22710 18420
rect 19904 18312 21128 18340
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19521 18235 19579 18241
rect 19628 18244 19809 18272
rect 14323 18176 15148 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 8113 18139 8171 18145
rect 8113 18136 8125 18139
rect 6472 18108 8125 18136
rect 8113 18105 8125 18108
rect 8159 18105 8171 18139
rect 8113 18099 8171 18105
rect 4154 18068 4160 18080
rect 3160 18040 4160 18068
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 5626 18028 5632 18080
rect 5684 18028 5690 18080
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 7156 18040 7205 18068
rect 7156 18028 7162 18040
rect 7193 18037 7205 18040
rect 7239 18037 7251 18071
rect 7193 18031 7251 18037
rect 8386 18028 8392 18080
rect 8444 18028 8450 18080
rect 11974 18028 11980 18080
rect 12032 18028 12038 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 14752 18068 14780 18176
rect 15286 18164 15292 18216
rect 15344 18164 15350 18216
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 15436 18176 15485 18204
rect 15436 18164 15442 18176
rect 15473 18173 15485 18176
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 16114 18164 16120 18216
rect 16172 18164 16178 18216
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 18506 18204 18512 18216
rect 17788 18176 18512 18204
rect 14829 18139 14887 18145
rect 14829 18105 14841 18139
rect 14875 18136 14887 18139
rect 14918 18136 14924 18148
rect 14875 18108 14924 18136
rect 14875 18105 14887 18108
rect 14829 18099 14887 18105
rect 14918 18096 14924 18108
rect 14976 18096 14982 18148
rect 17310 18096 17316 18148
rect 17368 18136 17374 18148
rect 17788 18136 17816 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 18690 18213 18696 18216
rect 18668 18207 18696 18213
rect 18668 18173 18680 18207
rect 18668 18167 18696 18173
rect 18690 18164 18696 18167
rect 18748 18164 18754 18216
rect 17368 18108 17816 18136
rect 19061 18139 19119 18145
rect 17368 18096 17374 18108
rect 19061 18105 19073 18139
rect 19107 18136 19119 18139
rect 19150 18136 19156 18148
rect 19107 18108 19156 18136
rect 19107 18105 19119 18108
rect 19061 18099 19119 18105
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 12492 18040 14780 18068
rect 17865 18071 17923 18077
rect 12492 18028 12498 18040
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 19628 18068 19656 18244
rect 19797 18241 19809 18244
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 20073 18275 20131 18281
rect 20073 18241 20085 18275
rect 20119 18272 20131 18275
rect 20162 18272 20168 18284
rect 20119 18244 20168 18272
rect 20119 18241 20131 18244
rect 20073 18235 20131 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20346 18281 20352 18284
rect 20340 18235 20352 18281
rect 20346 18232 20352 18235
rect 20404 18232 20410 18284
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 19886 18204 19892 18216
rect 19751 18176 19892 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 21100 18204 21128 18312
rect 22646 18281 22652 18284
rect 22624 18275 22652 18281
rect 22624 18241 22636 18275
rect 22624 18235 22652 18241
rect 22646 18232 22652 18235
rect 22704 18232 22710 18284
rect 22465 18207 22523 18213
rect 22465 18204 22477 18207
rect 21100 18176 22477 18204
rect 22002 18096 22008 18148
rect 22060 18136 22066 18148
rect 22103 18136 22131 18176
rect 22465 18173 22477 18176
rect 22511 18173 22523 18207
rect 22465 18167 22523 18173
rect 22741 18207 22799 18213
rect 22741 18173 22753 18207
rect 22787 18204 22799 18207
rect 22922 18204 22928 18216
rect 22787 18176 22928 18204
rect 22787 18173 22799 18176
rect 22741 18167 22799 18173
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 23474 18164 23480 18216
rect 23532 18164 23538 18216
rect 23661 18207 23719 18213
rect 23661 18173 23673 18207
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 22060 18108 22131 18136
rect 23017 18139 23075 18145
rect 22060 18096 22066 18108
rect 23017 18105 23029 18139
rect 23063 18105 23075 18139
rect 23017 18099 23075 18105
rect 17911 18040 19656 18068
rect 21821 18071 21879 18077
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 21821 18037 21833 18071
rect 21867 18068 21879 18071
rect 22554 18068 22560 18080
rect 21867 18040 22560 18068
rect 21867 18037 21879 18040
rect 21821 18031 21879 18037
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 22922 18028 22928 18080
rect 22980 18068 22986 18080
rect 23032 18068 23060 18099
rect 23106 18096 23112 18148
rect 23164 18136 23170 18148
rect 23676 18136 23704 18167
rect 23164 18108 23704 18136
rect 23164 18096 23170 18108
rect 22980 18040 23060 18068
rect 22980 18028 22986 18040
rect 1104 17978 24012 18000
rect 1104 17926 1350 17978
rect 1402 17926 1414 17978
rect 1466 17926 1478 17978
rect 1530 17926 1542 17978
rect 1594 17926 1606 17978
rect 1658 17926 4350 17978
rect 4402 17926 4414 17978
rect 4466 17926 4478 17978
rect 4530 17926 4542 17978
rect 4594 17926 4606 17978
rect 4658 17926 7350 17978
rect 7402 17926 7414 17978
rect 7466 17926 7478 17978
rect 7530 17926 7542 17978
rect 7594 17926 7606 17978
rect 7658 17926 10350 17978
rect 10402 17926 10414 17978
rect 10466 17926 10478 17978
rect 10530 17926 10542 17978
rect 10594 17926 10606 17978
rect 10658 17926 13350 17978
rect 13402 17926 13414 17978
rect 13466 17926 13478 17978
rect 13530 17926 13542 17978
rect 13594 17926 13606 17978
rect 13658 17926 16350 17978
rect 16402 17926 16414 17978
rect 16466 17926 16478 17978
rect 16530 17926 16542 17978
rect 16594 17926 16606 17978
rect 16658 17926 19350 17978
rect 19402 17926 19414 17978
rect 19466 17926 19478 17978
rect 19530 17926 19542 17978
rect 19594 17926 19606 17978
rect 19658 17926 22350 17978
rect 22402 17926 22414 17978
rect 22466 17926 22478 17978
rect 22530 17926 22542 17978
rect 22594 17926 22606 17978
rect 22658 17926 24012 17978
rect 1104 17904 24012 17926
rect 6733 17867 6791 17873
rect 6733 17833 6745 17867
rect 6779 17864 6791 17867
rect 6914 17864 6920 17876
rect 6779 17836 6920 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7285 17867 7343 17873
rect 7285 17833 7297 17867
rect 7331 17864 7343 17867
rect 7742 17864 7748 17876
rect 7331 17836 7748 17864
rect 7331 17833 7343 17836
rect 7285 17827 7343 17833
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 9125 17867 9183 17873
rect 9125 17833 9137 17867
rect 9171 17864 9183 17867
rect 11054 17864 11060 17876
rect 9171 17836 11060 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 14182 17864 14188 17876
rect 13495 17836 14188 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 14182 17824 14188 17836
rect 14240 17864 14246 17876
rect 14550 17864 14556 17876
rect 14240 17836 14556 17864
rect 14240 17824 14246 17836
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 15933 17867 15991 17873
rect 15933 17864 15945 17867
rect 15344 17836 15945 17864
rect 15344 17824 15350 17836
rect 15933 17833 15945 17836
rect 15979 17833 15991 17867
rect 15933 17827 15991 17833
rect 17678 17824 17684 17876
rect 17736 17864 17742 17876
rect 17773 17867 17831 17873
rect 17773 17864 17785 17867
rect 17736 17836 17785 17864
rect 17736 17824 17742 17836
rect 17773 17833 17785 17836
rect 17819 17833 17831 17867
rect 17773 17827 17831 17833
rect 19245 17867 19303 17873
rect 19245 17833 19257 17867
rect 19291 17864 19303 17867
rect 19702 17864 19708 17876
rect 19291 17836 19708 17864
rect 19291 17833 19303 17836
rect 19245 17827 19303 17833
rect 19702 17824 19708 17836
rect 19760 17824 19766 17876
rect 23106 17824 23112 17876
rect 23164 17824 23170 17876
rect 8757 17799 8815 17805
rect 8757 17765 8769 17799
rect 8803 17765 8815 17799
rect 8757 17759 8815 17765
rect 8772 17728 8800 17759
rect 17494 17756 17500 17808
rect 17552 17796 17558 17808
rect 17552 17768 18368 17796
rect 17552 17756 17558 17768
rect 9582 17728 9588 17740
rect 8772 17700 9588 17728
rect 9582 17688 9588 17700
rect 9640 17728 9646 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9640 17700 10057 17728
rect 9640 17688 9646 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10226 17688 10232 17740
rect 10284 17728 10290 17740
rect 10321 17731 10379 17737
rect 10321 17728 10333 17731
rect 10284 17700 10333 17728
rect 10284 17688 10290 17700
rect 10321 17697 10333 17700
rect 10367 17728 10379 17731
rect 10686 17728 10692 17740
rect 10367 17700 10692 17728
rect 10367 17697 10379 17700
rect 10321 17691 10379 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17728 10839 17731
rect 10870 17728 10876 17740
rect 10827 17700 10876 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11480 17700 11621 17728
rect 11480 17688 11486 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11756 17700 12081 17728
rect 11756 17688 11762 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 4212 17632 5365 17660
rect 4212 17620 4218 17632
rect 5353 17629 5365 17632
rect 5399 17660 5411 17663
rect 5399 17632 5764 17660
rect 5399 17629 5411 17632
rect 5353 17623 5411 17629
rect 5626 17601 5632 17604
rect 5620 17592 5632 17601
rect 5587 17564 5632 17592
rect 5620 17555 5632 17564
rect 5626 17552 5632 17555
rect 5684 17552 5690 17604
rect 5736 17592 5764 17632
rect 7098 17620 7104 17672
rect 7156 17620 7162 17672
rect 7190 17620 7196 17672
rect 7248 17660 7254 17672
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 7248 17632 7389 17660
rect 7248 17620 7254 17632
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 9858 17620 9864 17672
rect 9916 17669 9922 17672
rect 9916 17663 9965 17669
rect 9916 17629 9919 17663
rect 9953 17629 9965 17663
rect 9916 17623 9965 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11330 17660 11336 17672
rect 11011 17632 11336 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 9916 17620 9922 17623
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11974 17620 11980 17672
rect 12032 17660 12038 17672
rect 12325 17663 12383 17669
rect 12325 17660 12337 17663
rect 12032 17632 12337 17660
rect 12032 17620 12038 17632
rect 12325 17629 12337 17632
rect 12371 17629 12383 17663
rect 12325 17623 12383 17629
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17660 13783 17663
rect 14090 17660 14096 17672
rect 13771 17632 14096 17660
rect 13771 17629 13783 17632
rect 13725 17623 13783 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14182 17620 14188 17672
rect 14240 17620 14246 17672
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17660 14611 17663
rect 14642 17660 14648 17672
rect 14599 17632 14648 17660
rect 14599 17629 14611 17632
rect 14553 17623 14611 17629
rect 14642 17620 14648 17632
rect 14700 17660 14706 17672
rect 16301 17663 16359 17669
rect 16301 17660 16313 17663
rect 14700 17632 16313 17660
rect 14700 17620 14706 17632
rect 16301 17629 16313 17632
rect 16347 17660 16359 17663
rect 17402 17660 17408 17672
rect 16347 17632 17408 17660
rect 16347 17629 16359 17632
rect 16301 17623 16359 17629
rect 17402 17620 17408 17632
rect 17460 17620 17466 17672
rect 7208 17592 7236 17620
rect 5736 17564 7236 17592
rect 7644 17595 7702 17601
rect 7644 17561 7656 17595
rect 7690 17592 7702 17595
rect 7742 17592 7748 17604
rect 7690 17564 7748 17592
rect 7690 17561 7702 17564
rect 7644 17555 7702 17561
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 14826 17601 14832 17604
rect 11425 17595 11483 17601
rect 11425 17592 11437 17595
rect 10796 17564 11437 17592
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 10796 17524 10824 17564
rect 11425 17561 11437 17564
rect 11471 17561 11483 17595
rect 14820 17592 14832 17601
rect 14787 17564 14832 17592
rect 11425 17555 11483 17561
rect 14820 17555 14832 17564
rect 14826 17552 14832 17555
rect 14884 17552 14890 17604
rect 16568 17595 16626 17601
rect 16568 17561 16580 17595
rect 16614 17592 16626 17595
rect 16942 17592 16948 17604
rect 16614 17564 16948 17592
rect 16614 17561 16626 17564
rect 16568 17555 16626 17561
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 8720 17496 10824 17524
rect 8720 17484 8726 17496
rect 11054 17484 11060 17536
rect 11112 17484 11118 17536
rect 11514 17484 11520 17536
rect 11572 17484 11578 17536
rect 13538 17484 13544 17536
rect 13596 17484 13602 17536
rect 13814 17484 13820 17536
rect 13872 17524 13878 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 13872 17496 14381 17524
rect 13872 17484 13878 17496
rect 14369 17493 14381 17496
rect 14415 17524 14427 17527
rect 17512 17524 17540 17756
rect 18230 17688 18236 17740
rect 18288 17688 18294 17740
rect 18340 17737 18368 17768
rect 21192 17768 21772 17796
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17697 18383 17731
rect 19242 17728 19248 17740
rect 18325 17691 18383 17697
rect 18708 17700 19248 17728
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 17736 17632 18153 17660
rect 17736 17620 17742 17632
rect 18141 17629 18153 17632
rect 18187 17660 18199 17663
rect 18506 17660 18512 17672
rect 18187 17632 18512 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18506 17620 18512 17632
rect 18564 17660 18570 17672
rect 18708 17660 18736 17700
rect 19242 17688 19248 17700
rect 19300 17688 19306 17740
rect 21192 17737 21220 17768
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 21361 17731 21419 17737
rect 21361 17697 21373 17731
rect 21407 17728 21419 17731
rect 21634 17728 21640 17740
rect 21407 17700 21640 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 21744 17728 21772 17768
rect 21744 17700 21864 17728
rect 18564 17632 18736 17660
rect 18564 17620 18570 17632
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 20622 17660 20628 17672
rect 20180 17632 20628 17660
rect 20180 17604 20208 17632
rect 20622 17620 20628 17632
rect 20680 17660 20686 17672
rect 21729 17663 21787 17669
rect 21729 17660 21741 17663
rect 20680 17632 21741 17660
rect 20680 17620 20686 17632
rect 21729 17629 21741 17632
rect 21775 17629 21787 17663
rect 21836 17660 21864 17700
rect 21836 17632 22094 17660
rect 21729 17623 21787 17629
rect 18690 17592 18696 17604
rect 17696 17564 18696 17592
rect 17696 17533 17724 17564
rect 18690 17552 18696 17564
rect 18748 17552 18754 17604
rect 20162 17552 20168 17604
rect 20220 17552 20226 17604
rect 20254 17552 20260 17604
rect 20312 17592 20318 17604
rect 20358 17595 20416 17601
rect 20358 17592 20370 17595
rect 20312 17564 20370 17592
rect 20312 17552 20318 17564
rect 20358 17561 20370 17564
rect 20404 17561 20416 17595
rect 20358 17555 20416 17561
rect 21085 17595 21143 17601
rect 21085 17561 21097 17595
rect 21131 17592 21143 17595
rect 21131 17564 21588 17592
rect 21131 17561 21143 17564
rect 21085 17555 21143 17561
rect 14415 17496 17540 17524
rect 17681 17527 17739 17533
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 17681 17493 17693 17527
rect 17727 17493 17739 17527
rect 17681 17487 17739 17493
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 20530 17484 20536 17536
rect 20588 17524 20594 17536
rect 20717 17527 20775 17533
rect 20717 17524 20729 17527
rect 20588 17496 20729 17524
rect 20588 17484 20594 17496
rect 20717 17493 20729 17496
rect 20763 17493 20775 17527
rect 21560 17524 21588 17564
rect 21818 17552 21824 17604
rect 21876 17592 21882 17604
rect 21974 17595 22032 17601
rect 21974 17592 21986 17595
rect 21876 17564 21986 17592
rect 21876 17552 21882 17564
rect 21974 17561 21986 17564
rect 22020 17561 22032 17595
rect 22066 17592 22094 17632
rect 22278 17620 22284 17672
rect 22336 17660 22342 17672
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 22336 17632 23397 17660
rect 22336 17620 22342 17632
rect 23385 17629 23397 17632
rect 23431 17629 23443 17663
rect 23385 17623 23443 17629
rect 22738 17592 22744 17604
rect 22066 17564 22744 17592
rect 21974 17555 22032 17561
rect 22738 17552 22744 17564
rect 22796 17552 22802 17604
rect 22094 17524 22100 17536
rect 21560 17496 22100 17524
rect 20717 17487 20775 17493
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 23382 17484 23388 17536
rect 23440 17524 23446 17536
rect 23569 17527 23627 17533
rect 23569 17524 23581 17527
rect 23440 17496 23581 17524
rect 23440 17484 23446 17496
rect 23569 17493 23581 17496
rect 23615 17493 23627 17527
rect 23569 17487 23627 17493
rect 1104 17434 24164 17456
rect 1104 17382 2850 17434
rect 2902 17382 2914 17434
rect 2966 17382 2978 17434
rect 3030 17382 3042 17434
rect 3094 17382 3106 17434
rect 3158 17382 5850 17434
rect 5902 17382 5914 17434
rect 5966 17382 5978 17434
rect 6030 17382 6042 17434
rect 6094 17382 6106 17434
rect 6158 17382 8850 17434
rect 8902 17382 8914 17434
rect 8966 17382 8978 17434
rect 9030 17382 9042 17434
rect 9094 17382 9106 17434
rect 9158 17382 11850 17434
rect 11902 17382 11914 17434
rect 11966 17382 11978 17434
rect 12030 17382 12042 17434
rect 12094 17382 12106 17434
rect 12158 17382 14850 17434
rect 14902 17382 14914 17434
rect 14966 17382 14978 17434
rect 15030 17382 15042 17434
rect 15094 17382 15106 17434
rect 15158 17382 17850 17434
rect 17902 17382 17914 17434
rect 17966 17382 17978 17434
rect 18030 17382 18042 17434
rect 18094 17382 18106 17434
rect 18158 17382 20850 17434
rect 20902 17382 20914 17434
rect 20966 17382 20978 17434
rect 21030 17382 21042 17434
rect 21094 17382 21106 17434
rect 21158 17382 23850 17434
rect 23902 17382 23914 17434
rect 23966 17382 23978 17434
rect 24030 17382 24042 17434
rect 24094 17382 24106 17434
rect 24158 17382 24164 17434
rect 1104 17360 24164 17382
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5718 17320 5724 17332
rect 5316 17292 5724 17320
rect 5316 17280 5322 17292
rect 5718 17280 5724 17292
rect 5776 17320 5782 17332
rect 6822 17320 6828 17332
rect 5776 17292 6828 17320
rect 5776 17280 5782 17292
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 8662 17280 8668 17332
rect 8720 17280 8726 17332
rect 10778 17320 10784 17332
rect 8772 17292 10784 17320
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 8772 17252 8800 17292
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11330 17280 11336 17332
rect 11388 17280 11394 17332
rect 11514 17280 11520 17332
rect 11572 17280 11578 17332
rect 14645 17323 14703 17329
rect 14645 17289 14657 17323
rect 14691 17320 14703 17323
rect 15378 17320 15384 17332
rect 14691 17292 15384 17320
rect 14691 17289 14703 17292
rect 14645 17283 14703 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 16761 17323 16819 17329
rect 16761 17289 16773 17323
rect 16807 17320 16819 17323
rect 16850 17320 16856 17332
rect 16807 17292 16856 17320
rect 16807 17289 16819 17292
rect 16761 17283 16819 17289
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 17221 17323 17279 17329
rect 17221 17289 17233 17323
rect 17267 17289 17279 17323
rect 17221 17283 17279 17289
rect 17589 17323 17647 17329
rect 17589 17289 17601 17323
rect 17635 17320 17647 17323
rect 17770 17320 17776 17332
rect 17635 17292 17776 17320
rect 17635 17289 17647 17292
rect 17589 17283 17647 17289
rect 6604 17224 8800 17252
rect 6604 17212 6610 17224
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 9732 17224 9996 17252
rect 9732 17212 9738 17224
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17184 5319 17187
rect 5534 17184 5540 17196
rect 5307 17156 5540 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 5626 17144 5632 17196
rect 5684 17184 5690 17196
rect 9968 17193 9996 17224
rect 10226 17193 10232 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5684 17156 5733 17184
rect 5684 17144 5690 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 5859 17156 6377 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8757 17187 8815 17193
rect 8251 17156 8524 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17085 6055 17119
rect 5997 17079 6055 17085
rect 4246 17008 4252 17060
rect 4304 17048 4310 17060
rect 5718 17048 5724 17060
rect 4304 17020 5724 17048
rect 4304 17008 4310 17020
rect 5718 17008 5724 17020
rect 5776 17008 5782 17060
rect 6012 17048 6040 17079
rect 6454 17076 6460 17128
rect 6512 17116 6518 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6512 17088 6929 17116
rect 6512 17076 6518 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 7944 17116 7972 17147
rect 8386 17116 8392 17128
rect 7944 17088 8392 17116
rect 6917 17079 6975 17085
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 6546 17048 6552 17060
rect 6012 17020 6552 17048
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 6730 17008 6736 17060
rect 6788 17048 6794 17060
rect 8297 17051 8355 17057
rect 6788 17020 8156 17048
rect 6788 17008 6794 17020
rect 5074 16940 5080 16992
rect 5132 16940 5138 16992
rect 5353 16983 5411 16989
rect 5353 16949 5365 16983
rect 5399 16980 5411 16983
rect 5442 16980 5448 16992
rect 5399 16952 5448 16980
rect 5399 16949 5411 16952
rect 5353 16943 5411 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 8018 16940 8024 16992
rect 8076 16940 8082 16992
rect 8128 16980 8156 17020
rect 8297 17017 8309 17051
rect 8343 17048 8355 17051
rect 8496 17048 8524 17156
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8803 17156 9137 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10220 17147 10232 17193
rect 10226 17144 10232 17147
rect 10284 17144 10290 17196
rect 11348 17184 11376 17280
rect 11698 17212 11704 17264
rect 11756 17252 11762 17264
rect 12342 17252 12348 17264
rect 11756 17224 12348 17252
rect 11756 17212 11762 17224
rect 12342 17212 12348 17224
rect 12400 17252 12406 17264
rect 13538 17261 13544 17264
rect 13532 17252 13544 17261
rect 12400 17224 13308 17252
rect 13499 17224 13544 17252
rect 12400 17212 12406 17224
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11348 17156 12081 17184
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12710 17184 12716 17196
rect 12483 17156 12716 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13280 17193 13308 17224
rect 13532 17215 13544 17224
rect 13538 17212 13544 17215
rect 13596 17212 13602 17264
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 15378 17144 15384 17196
rect 15436 17144 15442 17196
rect 15470 17144 15476 17196
rect 15528 17144 15534 17196
rect 16945 17187 17003 17193
rect 16945 17153 16957 17187
rect 16991 17184 17003 17187
rect 17236 17184 17264 17283
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 19886 17320 19892 17332
rect 19475 17292 19892 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 20257 17323 20315 17329
rect 20257 17289 20269 17323
rect 20303 17320 20315 17323
rect 20346 17320 20352 17332
rect 20303 17292 20352 17320
rect 20303 17289 20315 17292
rect 20257 17283 20315 17289
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 22097 17323 22155 17329
rect 22097 17289 22109 17323
rect 22143 17320 22155 17323
rect 22278 17320 22284 17332
rect 22143 17292 22284 17320
rect 22143 17289 22155 17292
rect 22097 17283 22155 17289
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 23569 17323 23627 17329
rect 23569 17320 23581 17323
rect 23532 17292 23581 17320
rect 23532 17280 23538 17292
rect 23569 17289 23581 17292
rect 23615 17289 23627 17323
rect 23569 17283 23627 17289
rect 17402 17212 17408 17264
rect 17460 17252 17466 17264
rect 18316 17255 18374 17261
rect 17460 17224 18092 17252
rect 17460 17212 17466 17224
rect 16991 17156 17264 17184
rect 16991 17153 17003 17156
rect 16945 17147 17003 17153
rect 17678 17144 17684 17196
rect 17736 17144 17742 17196
rect 18064 17193 18092 17224
rect 18316 17221 18328 17255
rect 18362 17252 18374 17255
rect 18598 17252 18604 17264
rect 18362 17224 18604 17252
rect 18362 17221 18374 17224
rect 18316 17215 18374 17221
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 19904 17184 19932 17280
rect 20622 17212 20628 17264
rect 20680 17252 20686 17264
rect 21453 17255 21511 17261
rect 21453 17252 21465 17255
rect 20680 17224 21465 17252
rect 20680 17212 20686 17224
rect 21453 17221 21465 17224
rect 21499 17252 21511 17255
rect 22456 17255 22514 17261
rect 21499 17224 22094 17252
rect 21499 17221 21511 17224
rect 21453 17215 21511 17221
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 19904 17156 20085 17184
rect 18049 17147 18107 17153
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20441 17187 20499 17193
rect 20441 17153 20453 17187
rect 20487 17184 20499 17187
rect 20530 17184 20536 17196
rect 20487 17156 20536 17184
rect 20487 17153 20499 17156
rect 20441 17147 20499 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20714 17144 20720 17196
rect 20772 17144 20778 17196
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 21913 17187 21971 17193
rect 21913 17184 21925 17187
rect 21324 17156 21925 17184
rect 21324 17144 21330 17156
rect 21913 17153 21925 17156
rect 21959 17153 21971 17187
rect 22066 17184 22094 17224
rect 22456 17221 22468 17255
rect 22502 17252 22514 17255
rect 23198 17252 23204 17264
rect 22502 17224 23204 17252
rect 22502 17221 22514 17224
rect 22456 17215 22514 17221
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 22189 17187 22247 17193
rect 22189 17184 22201 17187
rect 22066 17156 22201 17184
rect 21913 17147 21971 17153
rect 22189 17153 22201 17156
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17116 8999 17119
rect 9490 17116 9496 17128
rect 8987 17088 9496 17116
rect 8987 17085 8999 17088
rect 8941 17079 8999 17085
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 9858 17116 9864 17128
rect 9732 17088 9864 17116
rect 9732 17076 9738 17088
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 17773 17119 17831 17125
rect 17773 17085 17785 17119
rect 17819 17085 17831 17119
rect 17773 17079 17831 17085
rect 8343 17020 8524 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 14550 17008 14556 17060
rect 14608 17048 14614 17060
rect 14737 17051 14795 17057
rect 14737 17048 14749 17051
rect 14608 17020 14749 17048
rect 14608 17008 14614 17020
rect 14737 17017 14749 17020
rect 14783 17017 14795 17051
rect 14737 17011 14795 17017
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 17788 17048 17816 17079
rect 15712 17020 17816 17048
rect 15712 17008 15718 17020
rect 19058 17008 19064 17060
rect 19116 17048 19122 17060
rect 19521 17051 19579 17057
rect 19521 17048 19533 17051
rect 19116 17020 19533 17048
rect 19116 17008 19122 17020
rect 19521 17017 19533 17020
rect 19567 17017 19579 17051
rect 19521 17011 19579 17017
rect 10134 16980 10140 16992
rect 8128 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 1104 16890 24012 16912
rect 1104 16838 1350 16890
rect 1402 16838 1414 16890
rect 1466 16838 1478 16890
rect 1530 16838 1542 16890
rect 1594 16838 1606 16890
rect 1658 16838 4350 16890
rect 4402 16838 4414 16890
rect 4466 16838 4478 16890
rect 4530 16838 4542 16890
rect 4594 16838 4606 16890
rect 4658 16838 7350 16890
rect 7402 16838 7414 16890
rect 7466 16838 7478 16890
rect 7530 16838 7542 16890
rect 7594 16838 7606 16890
rect 7658 16838 10350 16890
rect 10402 16838 10414 16890
rect 10466 16838 10478 16890
rect 10530 16838 10542 16890
rect 10594 16838 10606 16890
rect 10658 16838 13350 16890
rect 13402 16838 13414 16890
rect 13466 16838 13478 16890
rect 13530 16838 13542 16890
rect 13594 16838 13606 16890
rect 13658 16838 16350 16890
rect 16402 16838 16414 16890
rect 16466 16838 16478 16890
rect 16530 16838 16542 16890
rect 16594 16838 16606 16890
rect 16658 16838 19350 16890
rect 19402 16838 19414 16890
rect 19466 16838 19478 16890
rect 19530 16838 19542 16890
rect 19594 16838 19606 16890
rect 19658 16838 22350 16890
rect 22402 16838 22414 16890
rect 22466 16838 22478 16890
rect 22530 16838 22542 16890
rect 22594 16838 22606 16890
rect 22658 16838 24012 16890
rect 1104 16816 24012 16838
rect 4617 16779 4675 16785
rect 4617 16745 4629 16779
rect 4663 16776 4675 16779
rect 4663 16748 6776 16776
rect 4663 16745 4675 16748
rect 4617 16739 4675 16745
rect 5813 16711 5871 16717
rect 5813 16677 5825 16711
rect 5859 16708 5871 16711
rect 6638 16708 6644 16720
rect 5859 16680 6644 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 3973 16643 4031 16649
rect 3973 16640 3985 16643
rect 3936 16612 3985 16640
rect 3936 16600 3942 16612
rect 3973 16609 3985 16612
rect 4019 16640 4031 16643
rect 5399 16643 5457 16649
rect 5399 16640 5411 16643
rect 4019 16612 5411 16640
rect 4019 16609 4031 16612
rect 3973 16603 4031 16609
rect 5399 16609 5411 16612
rect 5445 16609 5457 16643
rect 5399 16603 5457 16609
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 5718 16640 5724 16652
rect 5583 16612 5724 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6454 16600 6460 16652
rect 6512 16600 6518 16652
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2774 16572 2780 16584
rect 2271 16544 2780 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 1302 16396 1308 16448
rect 1360 16436 1366 16448
rect 1489 16439 1547 16445
rect 1489 16436 1501 16439
rect 1360 16408 1501 16436
rect 1360 16396 1366 16408
rect 1489 16405 1501 16408
rect 1535 16405 1547 16439
rect 1688 16436 1716 16535
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 5258 16532 5264 16584
rect 5316 16532 5322 16584
rect 6270 16532 6276 16584
rect 6328 16532 6334 16584
rect 6748 16581 6776 16748
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 9677 16779 9735 16785
rect 9677 16776 9689 16779
rect 6880 16748 9689 16776
rect 6880 16736 6886 16748
rect 9677 16745 9689 16748
rect 9723 16776 9735 16779
rect 9766 16776 9772 16788
rect 9723 16748 9772 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 10226 16736 10232 16788
rect 10284 16736 10290 16788
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 11422 16776 11428 16788
rect 10836 16748 11428 16776
rect 10836 16736 10842 16748
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 14090 16736 14096 16788
rect 14148 16736 14154 16788
rect 18782 16736 18788 16788
rect 18840 16776 18846 16788
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 18840 16748 18981 16776
rect 18840 16736 18846 16748
rect 18969 16745 18981 16748
rect 19015 16745 19027 16779
rect 18969 16739 19027 16745
rect 20438 16736 20444 16788
rect 20496 16776 20502 16788
rect 20717 16779 20775 16785
rect 20717 16776 20729 16779
rect 20496 16748 20729 16776
rect 20496 16736 20502 16748
rect 20717 16745 20729 16748
rect 20763 16745 20775 16779
rect 20717 16739 20775 16745
rect 22094 16736 22100 16788
rect 22152 16736 22158 16788
rect 9217 16711 9275 16717
rect 9217 16677 9229 16711
rect 9263 16708 9275 16711
rect 9490 16708 9496 16720
rect 9263 16680 9496 16708
rect 9263 16677 9275 16680
rect 9217 16671 9275 16677
rect 9490 16668 9496 16680
rect 9548 16668 9554 16720
rect 22112 16708 22140 16736
rect 21376 16680 22508 16708
rect 7190 16600 7196 16652
rect 7248 16640 7254 16652
rect 7377 16643 7435 16649
rect 7377 16640 7389 16643
rect 7248 16612 7389 16640
rect 7248 16600 7254 16612
rect 7377 16609 7389 16612
rect 7423 16609 7435 16643
rect 11054 16640 11060 16652
rect 7377 16603 7435 16609
rect 10888 16612 11060 16640
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16541 6791 16575
rect 6733 16535 6791 16541
rect 7644 16575 7702 16581
rect 7644 16541 7656 16575
rect 7690 16572 7702 16575
rect 8018 16572 8024 16584
rect 7690 16544 8024 16572
rect 7690 16541 7702 16544
rect 7644 16535 7702 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16572 9459 16575
rect 9582 16572 9588 16584
rect 9447 16544 9588 16572
rect 9447 16541 9459 16544
rect 9401 16535 9459 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 10888 16572 10916 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 14550 16600 14556 16652
rect 14608 16600 14614 16652
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 18325 16643 18383 16649
rect 18325 16609 18337 16643
rect 18371 16609 18383 16643
rect 18325 16603 18383 16609
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16640 18567 16643
rect 19058 16640 19064 16652
rect 18555 16612 19064 16640
rect 18555 16609 18567 16612
rect 18509 16603 18567 16609
rect 10459 16544 10916 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 10962 16532 10968 16584
rect 11020 16572 11026 16584
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11020 16544 11805 16572
rect 11020 16532 11026 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 14366 16572 14372 16584
rect 11793 16535 11851 16541
rect 14292 16544 14372 16572
rect 2498 16513 2504 16516
rect 2492 16467 2504 16513
rect 2498 16464 2504 16467
rect 2556 16464 2562 16516
rect 9692 16504 9720 16532
rect 2746 16476 4752 16504
rect 2746 16436 2774 16476
rect 1688 16408 2774 16436
rect 3605 16439 3663 16445
rect 1489 16399 1547 16405
rect 3605 16405 3617 16439
rect 3651 16436 3663 16439
rect 4246 16436 4252 16448
rect 3651 16408 4252 16436
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 4246 16396 4252 16408
rect 4304 16396 4310 16448
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4488 16408 4537 16436
rect 4488 16396 4494 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4724 16436 4752 16476
rect 8772 16476 9720 16504
rect 9769 16507 9827 16513
rect 8772 16445 8800 16476
rect 9769 16473 9781 16507
rect 9815 16504 9827 16507
rect 12710 16504 12716 16516
rect 9815 16476 12716 16504
rect 9815 16473 9827 16476
rect 9769 16467 9827 16473
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 6549 16439 6607 16445
rect 6549 16436 6561 16439
rect 4724 16408 6561 16436
rect 4525 16399 4583 16405
rect 6549 16405 6561 16408
rect 6595 16405 6607 16439
rect 6549 16399 6607 16405
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16405 8815 16439
rect 8757 16399 8815 16405
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16436 11667 16439
rect 14292 16436 14320 16544
rect 14366 16532 14372 16544
rect 14424 16572 14430 16584
rect 14660 16572 14688 16603
rect 14424 16544 14688 16572
rect 16761 16575 16819 16581
rect 14424 16532 14430 16544
rect 16761 16541 16773 16575
rect 16807 16572 16819 16575
rect 16850 16572 16856 16584
rect 16807 16544 16856 16572
rect 16807 16541 16819 16544
rect 16761 16535 16819 16541
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 18340 16572 18368 16603
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 21232 16612 21281 16640
rect 21232 16600 21238 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 17736 16544 18368 16572
rect 17736 16532 17742 16544
rect 20622 16532 20628 16584
rect 20680 16532 20686 16584
rect 21082 16532 21088 16584
rect 21140 16532 21146 16584
rect 14458 16464 14464 16516
rect 14516 16464 14522 16516
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 18601 16507 18659 16513
rect 18601 16504 18613 16507
rect 18564 16476 18613 16504
rect 18564 16464 18570 16476
rect 18601 16473 18613 16476
rect 18647 16473 18659 16507
rect 18601 16467 18659 16473
rect 11655 16408 14320 16436
rect 11655 16405 11667 16408
rect 11609 16399 11667 16405
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 15988 16408 16129 16436
rect 15988 16396 15994 16408
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 16117 16399 16175 16405
rect 21177 16439 21235 16445
rect 21177 16405 21189 16439
rect 21223 16436 21235 16439
rect 21376 16436 21404 16680
rect 21726 16600 21732 16652
rect 21784 16640 21790 16652
rect 22186 16640 22192 16652
rect 21784 16612 22192 16640
rect 21784 16600 21790 16612
rect 22186 16600 22192 16612
rect 22244 16600 22250 16652
rect 21818 16532 21824 16584
rect 21876 16532 21882 16584
rect 22480 16581 22508 16680
rect 23474 16600 23480 16652
rect 23532 16600 23538 16652
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 22373 16507 22431 16513
rect 22373 16473 22385 16507
rect 22419 16504 22431 16507
rect 22925 16507 22983 16513
rect 22925 16504 22937 16507
rect 22419 16476 22937 16504
rect 22419 16473 22431 16476
rect 22373 16467 22431 16473
rect 22925 16473 22937 16476
rect 22971 16473 22983 16507
rect 22925 16467 22983 16473
rect 21223 16408 21404 16436
rect 22833 16439 22891 16445
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 22833 16405 22845 16439
rect 22879 16436 22891 16439
rect 23014 16436 23020 16448
rect 22879 16408 23020 16436
rect 22879 16405 22891 16408
rect 22833 16399 22891 16405
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 1104 16346 24164 16368
rect 1104 16294 2850 16346
rect 2902 16294 2914 16346
rect 2966 16294 2978 16346
rect 3030 16294 3042 16346
rect 3094 16294 3106 16346
rect 3158 16294 5850 16346
rect 5902 16294 5914 16346
rect 5966 16294 5978 16346
rect 6030 16294 6042 16346
rect 6094 16294 6106 16346
rect 6158 16294 8850 16346
rect 8902 16294 8914 16346
rect 8966 16294 8978 16346
rect 9030 16294 9042 16346
rect 9094 16294 9106 16346
rect 9158 16294 11850 16346
rect 11902 16294 11914 16346
rect 11966 16294 11978 16346
rect 12030 16294 12042 16346
rect 12094 16294 12106 16346
rect 12158 16294 14850 16346
rect 14902 16294 14914 16346
rect 14966 16294 14978 16346
rect 15030 16294 15042 16346
rect 15094 16294 15106 16346
rect 15158 16294 17850 16346
rect 17902 16294 17914 16346
rect 17966 16294 17978 16346
rect 18030 16294 18042 16346
rect 18094 16294 18106 16346
rect 18158 16294 20850 16346
rect 20902 16294 20914 16346
rect 20966 16294 20978 16346
rect 21030 16294 21042 16346
rect 21094 16294 21106 16346
rect 21158 16294 23850 16346
rect 23902 16294 23914 16346
rect 23966 16294 23978 16346
rect 24030 16294 24042 16346
rect 24094 16294 24106 16346
rect 24158 16294 24164 16346
rect 1104 16272 24164 16294
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2498 16232 2504 16244
rect 2455 16204 2504 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 2774 16232 2780 16244
rect 2746 16192 2780 16232
rect 2832 16192 2838 16244
rect 3878 16192 3884 16244
rect 3936 16192 3942 16244
rect 4430 16192 4436 16244
rect 4488 16192 4494 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6454 16232 6460 16244
rect 6227 16204 6460 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 15930 16192 15936 16244
rect 15988 16192 15994 16244
rect 20622 16192 20628 16244
rect 20680 16232 20686 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 20680 16204 23213 16232
rect 20680 16192 20686 16204
rect 23201 16201 23213 16204
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 2746 16164 2774 16192
rect 2516 16136 2774 16164
rect 750 16056 756 16108
rect 808 16096 814 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 808 16068 1409 16096
rect 808 16056 814 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 2222 16056 2228 16108
rect 2280 16056 2286 16108
rect 2516 16105 2544 16136
rect 2866 16124 2872 16176
rect 2924 16124 2930 16176
rect 5068 16167 5126 16173
rect 5068 16133 5080 16167
rect 5114 16164 5126 16167
rect 5258 16164 5264 16176
rect 5114 16136 5264 16164
rect 5114 16133 5126 16136
rect 5068 16127 5126 16133
rect 5258 16124 5264 16136
rect 5316 16124 5322 16176
rect 6270 16124 6276 16176
rect 6328 16164 6334 16176
rect 15841 16167 15899 16173
rect 6328 16136 7788 16164
rect 6328 16124 6334 16136
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16065 2559 16099
rect 2501 16059 2559 16065
rect 2768 16099 2826 16105
rect 2768 16065 2780 16099
rect 2814 16096 2826 16099
rect 2884 16096 2912 16124
rect 2814 16068 2912 16096
rect 4341 16099 4399 16105
rect 2814 16065 2826 16068
rect 2768 16059 2826 16065
rect 4341 16065 4353 16099
rect 4387 16096 4399 16099
rect 5626 16096 5632 16108
rect 4387 16068 5632 16096
rect 4387 16065 4399 16068
rect 4341 16059 4399 16065
rect 3510 15920 3516 15972
rect 3568 15960 3574 15972
rect 3973 15963 4031 15969
rect 3973 15960 3985 15963
rect 3568 15932 3985 15960
rect 3568 15920 3574 15932
rect 3973 15929 3985 15932
rect 4019 15929 4031 15963
rect 3973 15923 4031 15929
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 4154 15892 4160 15904
rect 1627 15864 4160 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 4154 15852 4160 15864
rect 4212 15892 4218 15904
rect 4356 15892 4384 16059
rect 5626 16056 5632 16068
rect 5684 16096 5690 16108
rect 7760 16105 7788 16136
rect 15841 16133 15853 16167
rect 15887 16164 15899 16167
rect 16022 16164 16028 16176
rect 15887 16136 16028 16164
rect 15887 16133 15899 16136
rect 15841 16127 15899 16133
rect 16022 16124 16028 16136
rect 16080 16164 16086 16176
rect 17589 16167 17647 16173
rect 17589 16164 17601 16167
rect 16080 16136 17601 16164
rect 16080 16124 16086 16136
rect 17589 16133 17601 16136
rect 17635 16164 17647 16167
rect 18782 16164 18788 16176
rect 17635 16136 18788 16164
rect 17635 16133 17647 16136
rect 17589 16127 17647 16133
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 20714 16124 20720 16176
rect 20772 16164 20778 16176
rect 21821 16167 21879 16173
rect 21821 16164 21833 16167
rect 20772 16136 21833 16164
rect 20772 16124 20778 16136
rect 21821 16133 21833 16136
rect 21867 16133 21879 16167
rect 21821 16127 21879 16133
rect 22186 16124 22192 16176
rect 22244 16164 22250 16176
rect 22244 16136 23428 16164
rect 22244 16124 22250 16136
rect 6733 16099 6791 16105
rect 6733 16096 6745 16099
rect 5684 16068 6745 16096
rect 5684 16056 5690 16068
rect 6733 16065 6745 16068
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6871 16068 7205 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 8294 16096 8300 16108
rect 8251 16068 8300 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 8294 16056 8300 16068
rect 8352 16096 8358 16108
rect 11882 16096 11888 16108
rect 8352 16068 11888 16096
rect 8352 16056 8358 16068
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16096 13139 16099
rect 13998 16096 14004 16108
rect 13127 16068 14004 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15562 16096 15568 16108
rect 15427 16068 15568 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 16298 16056 16304 16108
rect 16356 16096 16362 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16356 16068 16865 16096
rect 16356 16056 16362 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 17727 16068 18061 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16096 20039 16099
rect 20441 16099 20499 16105
rect 20027 16068 20116 16096
rect 20027 16065 20039 16068
rect 19981 16059 20039 16065
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 4706 16028 4712 16040
rect 4663 16000 4712 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 4798 15988 4804 16040
rect 4856 15988 4862 16040
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 6696 16000 6929 16028
rect 6696 15988 6702 16000
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 12529 16031 12587 16037
rect 12529 15997 12541 16031
rect 12575 16028 12587 16031
rect 12986 16028 12992 16040
rect 12575 16000 12992 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 12986 15988 12992 16000
rect 13044 15988 13050 16040
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 16206 16028 16212 16040
rect 16163 16000 16212 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 17773 16031 17831 16037
rect 17773 15997 17785 16031
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 9950 15920 9956 15972
rect 10008 15960 10014 15972
rect 13262 15960 13268 15972
rect 10008 15932 13268 15960
rect 10008 15920 10014 15932
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 16758 15920 16764 15972
rect 16816 15960 16822 15972
rect 17221 15963 17279 15969
rect 17221 15960 17233 15963
rect 16816 15932 17233 15960
rect 16816 15920 16822 15932
rect 17221 15929 17233 15932
rect 17267 15929 17279 15963
rect 17221 15923 17279 15929
rect 17678 15920 17684 15972
rect 17736 15960 17742 15972
rect 17788 15960 17816 15991
rect 18598 15988 18604 16040
rect 18656 15988 18662 16040
rect 20088 15969 20116 16068
rect 20441 16065 20453 16099
rect 20487 16096 20499 16099
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20487 16068 20913 16096
rect 20487 16065 20499 16068
rect 20441 16059 20499 16065
rect 20901 16065 20913 16068
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 21082 16056 21088 16108
rect 21140 16096 21146 16108
rect 21140 16068 22968 16096
rect 21140 16056 21146 16068
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 17736 15932 17816 15960
rect 20073 15963 20131 15969
rect 17736 15920 17742 15932
rect 20073 15929 20085 15963
rect 20119 15929 20131 15963
rect 20073 15923 20131 15929
rect 4212 15864 4384 15892
rect 4212 15852 4218 15864
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 5592 15864 6377 15892
rect 5592 15852 5598 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 6365 15855 6423 15861
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 8021 15895 8079 15901
rect 8021 15892 8033 15895
rect 7984 15864 8033 15892
rect 7984 15852 7990 15864
rect 8021 15861 8033 15864
rect 8067 15861 8079 15895
rect 8021 15855 8079 15861
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10962 15892 10968 15904
rect 10735 15864 10968 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11756 15864 11897 15892
rect 11756 15852 11762 15864
rect 11885 15861 11897 15864
rect 11931 15861 11943 15895
rect 11885 15855 11943 15861
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12860 15864 12909 15892
rect 12860 15852 12866 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 15197 15895 15255 15901
rect 15197 15892 15209 15895
rect 15160 15864 15209 15892
rect 15160 15852 15166 15864
rect 15197 15861 15209 15864
rect 15243 15861 15255 15895
rect 15197 15855 15255 15861
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 15436 15864 15485 15892
rect 15436 15852 15442 15864
rect 15473 15861 15485 15864
rect 15519 15861 15531 15895
rect 15473 15855 15531 15861
rect 17037 15895 17095 15901
rect 17037 15861 17049 15895
rect 17083 15892 17095 15895
rect 18966 15892 18972 15904
rect 17083 15864 18972 15892
rect 17083 15861 17095 15864
rect 17037 15855 17095 15861
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 19794 15852 19800 15904
rect 19852 15852 19858 15904
rect 20548 15892 20576 15991
rect 20640 15960 20668 15991
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 21453 16031 21511 16037
rect 21453 16028 21465 16031
rect 20772 16000 21465 16028
rect 20772 15988 20778 16000
rect 21453 15997 21465 16000
rect 21499 16028 21511 16031
rect 21910 16028 21916 16040
rect 21499 16000 21916 16028
rect 21499 15997 21511 16000
rect 21453 15991 21511 15997
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22066 16000 22569 16028
rect 21174 15960 21180 15972
rect 20640 15932 21180 15960
rect 21174 15920 21180 15932
rect 21232 15960 21238 15972
rect 21358 15960 21364 15972
rect 21232 15932 21364 15960
rect 21232 15920 21238 15932
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 21818 15920 21824 15972
rect 21876 15960 21882 15972
rect 22066 15960 22094 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 21876 15932 22094 15960
rect 21876 15920 21882 15932
rect 20622 15892 20628 15904
rect 20548 15864 20628 15892
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 22833 15895 22891 15901
rect 22833 15892 22845 15895
rect 20864 15864 22845 15892
rect 20864 15852 20870 15864
rect 22833 15861 22845 15864
rect 22879 15861 22891 15895
rect 22940 15892 22968 16068
rect 23400 16037 23428 16136
rect 23293 16031 23351 16037
rect 23293 15997 23305 16031
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 23308 15960 23336 15991
rect 23308 15932 24072 15960
rect 23658 15892 23664 15904
rect 22940 15864 23664 15892
rect 22833 15855 22891 15861
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 1104 15802 24012 15824
rect 1104 15750 1350 15802
rect 1402 15750 1414 15802
rect 1466 15750 1478 15802
rect 1530 15750 1542 15802
rect 1594 15750 1606 15802
rect 1658 15750 4350 15802
rect 4402 15750 4414 15802
rect 4466 15750 4478 15802
rect 4530 15750 4542 15802
rect 4594 15750 4606 15802
rect 4658 15750 7350 15802
rect 7402 15750 7414 15802
rect 7466 15750 7478 15802
rect 7530 15750 7542 15802
rect 7594 15750 7606 15802
rect 7658 15750 10350 15802
rect 10402 15750 10414 15802
rect 10466 15750 10478 15802
rect 10530 15750 10542 15802
rect 10594 15750 10606 15802
rect 10658 15750 13350 15802
rect 13402 15750 13414 15802
rect 13466 15750 13478 15802
rect 13530 15750 13542 15802
rect 13594 15750 13606 15802
rect 13658 15750 16350 15802
rect 16402 15750 16414 15802
rect 16466 15750 16478 15802
rect 16530 15750 16542 15802
rect 16594 15750 16606 15802
rect 16658 15750 19350 15802
rect 19402 15750 19414 15802
rect 19466 15750 19478 15802
rect 19530 15750 19542 15802
rect 19594 15750 19606 15802
rect 19658 15750 22350 15802
rect 22402 15750 22414 15802
rect 22466 15750 22478 15802
rect 22530 15750 22542 15802
rect 22594 15750 22606 15802
rect 22658 15750 24012 15802
rect 1104 15728 24012 15750
rect 2866 15648 2872 15700
rect 2924 15648 2930 15700
rect 6181 15691 6239 15697
rect 4448 15660 5764 15688
rect 2222 15580 2228 15632
rect 2280 15620 2286 15632
rect 3789 15623 3847 15629
rect 3789 15620 3801 15623
rect 2280 15592 3801 15620
rect 2280 15580 2286 15592
rect 3789 15589 3801 15592
rect 3835 15589 3847 15623
rect 3789 15583 3847 15589
rect 4448 15564 4476 15660
rect 5736 15620 5764 15660
rect 6181 15657 6193 15691
rect 6227 15688 6239 15691
rect 6270 15688 6276 15700
rect 6227 15660 6276 15688
rect 6227 15657 6239 15660
rect 6181 15651 6239 15657
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 14090 15688 14096 15700
rect 9732 15660 14096 15688
rect 9732 15648 9738 15660
rect 7926 15620 7932 15632
rect 5736 15592 7932 15620
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 8110 15580 8116 15632
rect 8168 15620 8174 15632
rect 8389 15623 8447 15629
rect 8389 15620 8401 15623
rect 8168 15592 8401 15620
rect 8168 15580 8174 15592
rect 8389 15589 8401 15592
rect 8435 15589 8447 15623
rect 8389 15583 8447 15589
rect 9769 15623 9827 15629
rect 9769 15589 9781 15623
rect 9815 15620 9827 15623
rect 10134 15620 10140 15632
rect 9815 15592 10140 15620
rect 9815 15589 9827 15592
rect 9769 15583 9827 15589
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 2832 15524 3832 15552
rect 2832 15512 2838 15524
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3510 15484 3516 15496
rect 3099 15456 3516 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 3804 15484 3832 15524
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 4249 15555 4307 15561
rect 4249 15552 4261 15555
rect 4212 15524 4261 15552
rect 4212 15512 4218 15524
rect 4249 15521 4261 15524
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8352 15524 8953 15552
rect 8352 15512 8358 15524
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 10962 15512 10968 15564
rect 11020 15512 11026 15564
rect 11164 15561 11192 15660
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 17494 15688 17500 15700
rect 16868 15660 17500 15688
rect 11514 15580 11520 15632
rect 11572 15620 11578 15632
rect 16209 15623 16267 15629
rect 11572 15592 12388 15620
rect 11572 15580 11578 15592
rect 12360 15564 12388 15592
rect 16209 15589 16221 15623
rect 16255 15620 16267 15623
rect 16868 15620 16896 15660
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 18739 15660 20392 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 16255 15592 16896 15620
rect 16255 15589 16267 15592
rect 16209 15583 16267 15589
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 11882 15552 11888 15564
rect 11480 15524 11888 15552
rect 11480 15512 11486 15524
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12342 15512 12348 15564
rect 12400 15512 12406 15564
rect 16666 15512 16672 15564
rect 16724 15512 16730 15564
rect 16868 15552 16896 15592
rect 17770 15580 17776 15632
rect 17828 15620 17834 15632
rect 19242 15620 19248 15632
rect 17828 15592 19248 15620
rect 17828 15580 17834 15592
rect 19242 15580 19248 15592
rect 19300 15580 19306 15632
rect 20364 15620 20392 15660
rect 20714 15648 20720 15700
rect 20772 15648 20778 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 21266 15688 21272 15700
rect 21131 15660 21272 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 23290 15688 23296 15700
rect 21376 15660 23296 15688
rect 21376 15620 21404 15660
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 23661 15691 23719 15697
rect 23661 15657 23673 15691
rect 23707 15688 23719 15691
rect 24044 15688 24072 15932
rect 23707 15660 24072 15688
rect 23707 15657 23719 15660
rect 23661 15651 23719 15657
rect 20364 15592 21404 15620
rect 22278 15580 22284 15632
rect 22336 15620 22342 15632
rect 22830 15620 22836 15632
rect 22336 15592 22836 15620
rect 22336 15580 22342 15592
rect 22830 15580 22836 15592
rect 22888 15580 22894 15632
rect 17034 15552 17040 15564
rect 16868 15524 17040 15552
rect 17034 15512 17040 15524
rect 17092 15512 17098 15564
rect 17209 15512 17215 15564
rect 17267 15552 17273 15564
rect 17267 15524 17311 15552
rect 17267 15512 17273 15524
rect 17494 15512 17500 15564
rect 17552 15512 17558 15564
rect 18417 15555 18475 15561
rect 18417 15521 18429 15555
rect 18463 15552 18475 15555
rect 18598 15552 18604 15564
rect 18463 15524 18604 15552
rect 18463 15521 18475 15524
rect 18417 15515 18475 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15552 21787 15555
rect 22186 15552 22192 15564
rect 21775 15524 22192 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 22186 15512 22192 15524
rect 22244 15512 22250 15564
rect 22741 15555 22799 15561
rect 22741 15521 22753 15555
rect 22787 15552 22799 15555
rect 22787 15524 23152 15552
rect 22787 15521 22799 15524
rect 22741 15515 22799 15521
rect 4798 15484 4804 15496
rect 3804 15456 4804 15484
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 5074 15493 5080 15496
rect 5068 15484 5080 15493
rect 5035 15456 5080 15484
rect 5068 15447 5080 15456
rect 5074 15444 5080 15447
rect 5132 15444 5138 15496
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 7742 15484 7748 15496
rect 7699 15456 7748 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 9674 15484 9680 15496
rect 8619 15456 9680 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 9950 15444 9956 15496
rect 10008 15444 10014 15496
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15102 15493 15108 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 14792 15456 14841 15484
rect 14792 15444 14798 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 15096 15484 15108 15493
rect 15063 15456 15108 15484
rect 14829 15447 14887 15453
rect 15096 15447 15108 15456
rect 15102 15444 15108 15447
rect 15160 15444 15166 15496
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15484 16359 15487
rect 16684 15484 16712 15512
rect 17402 15500 17408 15512
rect 17395 15493 17408 15500
rect 16347 15456 16712 15484
rect 17380 15487 17408 15493
rect 16347 15453 16359 15456
rect 16301 15447 16359 15453
rect 17380 15453 17392 15487
rect 17460 15460 17466 15512
rect 23124 15496 23152 15524
rect 17426 15453 17438 15460
rect 17380 15447 17438 15453
rect 18230 15444 18236 15496
rect 18288 15444 18294 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 7006 15416 7012 15428
rect 1596 15388 7012 15416
rect 1596 15357 1624 15388
rect 7006 15376 7012 15388
rect 7064 15416 7070 15428
rect 7558 15416 7564 15428
rect 7064 15388 7564 15416
rect 7064 15376 7070 15388
rect 7558 15376 7564 15388
rect 7616 15376 7622 15428
rect 10873 15419 10931 15425
rect 10873 15385 10885 15419
rect 10919 15416 10931 15419
rect 11793 15419 11851 15425
rect 11793 15416 11805 15419
rect 10919 15388 11805 15416
rect 10919 15385 10931 15388
rect 10873 15379 10931 15385
rect 11793 15385 11805 15388
rect 11839 15385 11851 15419
rect 11793 15379 11851 15385
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 8110 15348 8116 15360
rect 4764 15320 8116 15348
rect 4764 15308 4770 15320
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 8202 15308 8208 15360
rect 8260 15308 8266 15360
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10284 15320 10517 15348
rect 10284 15308 10290 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 10505 15311 10563 15317
rect 11330 15308 11336 15360
rect 11388 15308 11394 15360
rect 11808 15348 11836 15379
rect 12434 15376 12440 15428
rect 12492 15416 12498 15428
rect 12590 15419 12648 15425
rect 12590 15416 12602 15419
rect 12492 15388 12602 15416
rect 12492 15376 12498 15388
rect 12590 15385 12602 15388
rect 12636 15385 12648 15419
rect 12590 15379 12648 15385
rect 12894 15348 12900 15360
rect 11808 15320 12900 15348
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15348 13783 15351
rect 13906 15348 13912 15360
rect 13771 15320 13912 15348
rect 13771 15317 13783 15320
rect 13725 15311 13783 15317
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 16482 15308 16488 15360
rect 16540 15308 16546 15360
rect 16577 15351 16635 15357
rect 16577 15317 16589 15351
rect 16623 15348 16635 15351
rect 18524 15348 18552 15447
rect 19334 15444 19340 15496
rect 19392 15444 19398 15496
rect 20806 15444 20812 15496
rect 20864 15444 20870 15496
rect 21910 15493 21916 15496
rect 21888 15487 21916 15493
rect 21888 15453 21900 15487
rect 21888 15447 21916 15453
rect 21910 15444 21916 15447
rect 21968 15444 21974 15496
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15484 22983 15487
rect 23014 15484 23020 15496
rect 22971 15456 23020 15484
rect 22971 15453 22983 15456
rect 22925 15447 22983 15453
rect 23014 15444 23020 15456
rect 23072 15444 23078 15496
rect 23106 15444 23112 15496
rect 23164 15444 23170 15496
rect 19604 15419 19662 15425
rect 19604 15385 19616 15419
rect 19650 15416 19662 15419
rect 19794 15416 19800 15428
rect 19650 15388 19800 15416
rect 19650 15385 19662 15388
rect 19604 15379 19662 15385
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 21082 15416 21088 15428
rect 19904 15388 21088 15416
rect 16623 15320 18552 15348
rect 16623 15317 16635 15320
rect 16577 15311 16635 15317
rect 18782 15308 18788 15360
rect 18840 15348 18846 15360
rect 19904 15348 19932 15388
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 18840 15320 19932 15348
rect 20993 15351 21051 15357
rect 18840 15308 18846 15320
rect 20993 15317 21005 15351
rect 21039 15348 21051 15351
rect 21450 15348 21456 15360
rect 21039 15320 21456 15348
rect 21039 15317 21051 15320
rect 20993 15311 21051 15317
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 1104 15258 24164 15280
rect 1104 15206 2850 15258
rect 2902 15206 2914 15258
rect 2966 15206 2978 15258
rect 3030 15206 3042 15258
rect 3094 15206 3106 15258
rect 3158 15206 5850 15258
rect 5902 15206 5914 15258
rect 5966 15206 5978 15258
rect 6030 15206 6042 15258
rect 6094 15206 6106 15258
rect 6158 15206 8850 15258
rect 8902 15206 8914 15258
rect 8966 15206 8978 15258
rect 9030 15206 9042 15258
rect 9094 15206 9106 15258
rect 9158 15206 11850 15258
rect 11902 15206 11914 15258
rect 11966 15206 11978 15258
rect 12030 15206 12042 15258
rect 12094 15206 12106 15258
rect 12158 15206 14850 15258
rect 14902 15206 14914 15258
rect 14966 15206 14978 15258
rect 15030 15206 15042 15258
rect 15094 15206 15106 15258
rect 15158 15206 17850 15258
rect 17902 15206 17914 15258
rect 17966 15206 17978 15258
rect 18030 15206 18042 15258
rect 18094 15206 18106 15258
rect 18158 15206 20850 15258
rect 20902 15206 20914 15258
rect 20966 15206 20978 15258
rect 21030 15206 21042 15258
rect 21094 15206 21106 15258
rect 21158 15206 23850 15258
rect 23902 15206 23914 15258
rect 23966 15206 23978 15258
rect 24030 15206 24042 15258
rect 24094 15206 24106 15258
rect 24158 15206 24164 15258
rect 1104 15184 24164 15206
rect 3973 15147 4031 15153
rect 3973 15113 3985 15147
rect 4019 15144 4031 15147
rect 4154 15144 4160 15156
rect 4019 15116 4160 15144
rect 4019 15113 4031 15116
rect 3973 15107 4031 15113
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 5258 15104 5264 15156
rect 5316 15104 5322 15156
rect 7285 15147 7343 15153
rect 7285 15113 7297 15147
rect 7331 15113 7343 15147
rect 7285 15107 7343 15113
rect 4246 15036 4252 15088
rect 4304 15076 4310 15088
rect 4304 15048 4568 15076
rect 4304 15036 4310 15048
rect 1210 14968 1216 15020
rect 1268 15008 1274 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 1268 14980 1409 15008
rect 1268 14968 1274 14980
rect 1397 14977 1409 14980
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 2958 14968 2964 15020
rect 3016 15008 3022 15020
rect 3326 15008 3332 15020
rect 3016 14980 3332 15008
rect 3016 14968 3022 14980
rect 3326 14968 3332 14980
rect 3384 15008 3390 15020
rect 4430 15008 4436 15020
rect 3384 14980 4436 15008
rect 3384 14968 3390 14980
rect 4430 14968 4436 14980
rect 4488 14968 4494 15020
rect 4540 15017 4568 15048
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 5442 14968 5448 15020
rect 5500 14968 5506 15020
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 15008 7067 15011
rect 7300 15008 7328 15107
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 7616 15116 7665 15144
rect 7616 15104 7622 15116
rect 7653 15113 7665 15116
rect 7699 15113 7711 15147
rect 7653 15107 7711 15113
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 8202 15144 8208 15156
rect 7791 15116 8208 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9490 15144 9496 15156
rect 9416 15116 9496 15144
rect 9416 15076 9444 15116
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11333 15147 11391 15153
rect 11333 15144 11345 15147
rect 11296 15116 11345 15144
rect 11296 15104 11302 15116
rect 11333 15113 11345 15116
rect 11379 15113 11391 15147
rect 11333 15107 11391 15113
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15144 12035 15147
rect 12434 15144 12440 15156
rect 12023 15116 12440 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12434 15104 12440 15116
rect 12492 15104 12498 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13078 15144 13084 15156
rect 12952 15116 13084 15144
rect 12952 15104 12958 15116
rect 13078 15104 13084 15116
rect 13136 15144 13142 15156
rect 13136 15116 13768 15144
rect 13136 15104 13142 15116
rect 11514 15076 11520 15088
rect 7055 14980 7328 15008
rect 7852 15048 9444 15076
rect 9508 15048 11520 15076
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 4246 14940 4252 14952
rect 3651 14912 4252 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 4890 14900 4896 14952
rect 4948 14940 4954 14952
rect 7852 14949 7880 15048
rect 9237 15011 9295 15017
rect 9237 14977 9249 15011
rect 9283 15008 9295 15011
rect 9398 15008 9404 15020
rect 9283 14980 9404 15008
rect 9283 14977 9295 14980
rect 9237 14971 9295 14977
rect 9398 14968 9404 14980
rect 9456 14968 9462 15020
rect 9508 15017 9536 15048
rect 9968 15017 9996 15048
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 13740 15076 13768 15116
rect 13998 15104 14004 15156
rect 14056 15104 14062 15156
rect 16114 15144 16120 15156
rect 14660 15116 16120 15144
rect 14369 15079 14427 15085
rect 14369 15076 14381 15079
rect 13740 15048 14381 15076
rect 14369 15045 14381 15048
rect 14415 15045 14427 15079
rect 14369 15039 14427 15045
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 4948 14912 7849 14940
rect 4948 14900 4954 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 6638 14832 6644 14884
rect 6696 14872 6702 14884
rect 8113 14875 8171 14881
rect 6696 14844 8064 14872
rect 6696 14832 6702 14844
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 2682 14804 2688 14816
rect 1627 14776 2688 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 2866 14764 2872 14816
rect 2924 14804 2930 14816
rect 2961 14807 3019 14813
rect 2961 14804 2973 14807
rect 2924 14776 2973 14804
rect 2924 14764 2930 14776
rect 2961 14773 2973 14776
rect 3007 14773 3019 14807
rect 2961 14767 3019 14773
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 8036 14804 8064 14844
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 8294 14872 8300 14884
rect 8159 14844 8300 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 8294 14832 8300 14844
rect 8352 14832 8358 14884
rect 9122 14804 9128 14816
rect 8036 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14804 9186 14816
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 9180 14776 9689 14804
rect 9180 14764 9186 14776
rect 9677 14773 9689 14776
rect 9723 14773 9735 14807
rect 9876 14804 9904 14971
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10209 15011 10267 15017
rect 10209 15008 10221 15011
rect 10100 14980 10221 15008
rect 10100 14968 10106 14980
rect 10209 14977 10221 14980
rect 10255 14977 10267 15011
rect 10209 14971 10267 14977
rect 11330 14968 11336 15020
rect 11388 15008 11394 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11388 14980 11713 15008
rect 11388 14968 11394 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 12710 14968 12716 15020
rect 12768 14968 12774 15020
rect 12986 14968 12992 15020
rect 13044 14968 13050 15020
rect 14660 14952 14688 15116
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15144 16267 15147
rect 16850 15144 16856 15156
rect 16255 15116 16856 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16850 15104 16856 15116
rect 16908 15144 16914 15156
rect 17402 15144 17408 15156
rect 16908 15116 17408 15144
rect 16908 15104 16914 15116
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18598 15144 18604 15156
rect 18371 15116 18604 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18782 15104 18788 15156
rect 18840 15104 18846 15156
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 20438 15144 20444 15156
rect 19024 15116 20444 15144
rect 19024 15104 19030 15116
rect 20438 15104 20444 15116
rect 20496 15144 20502 15156
rect 21726 15144 21732 15156
rect 20496 15116 21732 15144
rect 20496 15104 20502 15116
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 23382 15104 23388 15156
rect 23440 15144 23446 15156
rect 23569 15147 23627 15153
rect 23569 15144 23581 15147
rect 23440 15116 23581 15144
rect 23440 15104 23446 15116
rect 23569 15113 23581 15116
rect 23615 15113 23627 15147
rect 23569 15107 23627 15113
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 14792 15048 16252 15076
rect 14792 15036 14798 15048
rect 14844 15017 14872 15048
rect 15102 15017 15108 15020
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 15096 14971 15108 15017
rect 15102 14968 15108 14971
rect 15160 14968 15166 15020
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 12851 14943 12909 14949
rect 12851 14940 12863 14943
rect 11296 14912 12863 14940
rect 11296 14900 11302 14912
rect 12851 14909 12863 14912
rect 12897 14909 12909 14943
rect 12851 14903 12909 14909
rect 13262 14900 13268 14952
rect 13320 14900 13326 14952
rect 13722 14900 13728 14952
rect 13780 14900 13786 14952
rect 13906 14900 13912 14952
rect 13964 14900 13970 14952
rect 14458 14900 14464 14952
rect 14516 14900 14522 14952
rect 14642 14900 14648 14952
rect 14700 14900 14706 14952
rect 16224 14940 16252 15048
rect 16482 15036 16488 15088
rect 16540 15076 16546 15088
rect 17190 15079 17248 15085
rect 17190 15076 17202 15079
rect 16540 15048 17202 15076
rect 16540 15036 16546 15048
rect 17190 15045 17202 15048
rect 17236 15045 17248 15079
rect 17190 15039 17248 15045
rect 21818 15036 21824 15088
rect 21876 15076 21882 15088
rect 21876 15048 23244 15076
rect 21876 15036 21882 15048
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 19604 15011 19662 15017
rect 16715 14980 18460 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16942 14940 16948 14952
rect 16224 14912 16948 14940
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 18432 14881 18460 14980
rect 19604 14977 19616 15011
rect 19650 15008 19662 15011
rect 19978 15008 19984 15020
rect 19650 14980 19984 15008
rect 19650 14977 19662 14980
rect 19604 14971 19662 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20772 14980 21189 15008
rect 20772 14968 20778 14980
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 22922 14968 22928 15020
rect 22980 15017 22986 15020
rect 23216 15017 23244 15048
rect 22980 14971 22992 15017
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23201 14971 23259 14977
rect 22980 14968 22986 14971
rect 23290 14968 23296 15020
rect 23348 15008 23354 15020
rect 23385 15011 23443 15017
rect 23385 15008 23397 15011
rect 23348 14980 23397 15008
rect 23348 14968 23354 14980
rect 23385 14977 23397 14980
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 18874 14900 18880 14952
rect 18932 14900 18938 14952
rect 18966 14900 18972 14952
rect 19024 14900 19030 14952
rect 19334 14900 19340 14952
rect 19392 14900 19398 14952
rect 20990 14900 20996 14952
rect 21048 14940 21054 14952
rect 21269 14943 21327 14949
rect 21269 14940 21281 14943
rect 21048 14912 21281 14940
rect 21048 14900 21054 14912
rect 21269 14909 21281 14912
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 21453 14943 21511 14949
rect 21453 14909 21465 14943
rect 21499 14940 21511 14943
rect 21634 14940 21640 14952
rect 21499 14912 21640 14940
rect 21499 14909 21511 14912
rect 21453 14903 21511 14909
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 18417 14875 18475 14881
rect 18417 14841 18429 14875
rect 18463 14841 18475 14875
rect 18417 14835 18475 14841
rect 20717 14875 20775 14881
rect 20717 14841 20729 14875
rect 20763 14872 20775 14875
rect 21910 14872 21916 14884
rect 20763 14844 21916 14872
rect 20763 14841 20775 14844
rect 20717 14835 20775 14841
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 11054 14804 11060 14816
rect 9876 14776 11060 14804
rect 9677 14767 9735 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 11514 14764 11520 14816
rect 11572 14764 11578 14816
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 14274 14804 14280 14816
rect 12115 14776 14280 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 16853 14807 16911 14813
rect 16853 14773 16865 14807
rect 16899 14804 16911 14807
rect 17218 14804 17224 14816
rect 16899 14776 17224 14804
rect 16899 14773 16911 14776
rect 16853 14767 16911 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 20806 14764 20812 14816
rect 20864 14764 20870 14816
rect 21821 14807 21879 14813
rect 21821 14773 21833 14807
rect 21867 14804 21879 14807
rect 23014 14804 23020 14816
rect 21867 14776 23020 14804
rect 21867 14773 21879 14776
rect 21821 14767 21879 14773
rect 23014 14764 23020 14776
rect 23072 14764 23078 14816
rect 1104 14714 24012 14736
rect 1104 14662 1350 14714
rect 1402 14662 1414 14714
rect 1466 14662 1478 14714
rect 1530 14662 1542 14714
rect 1594 14662 1606 14714
rect 1658 14662 4350 14714
rect 4402 14662 4414 14714
rect 4466 14662 4478 14714
rect 4530 14662 4542 14714
rect 4594 14662 4606 14714
rect 4658 14662 7350 14714
rect 7402 14662 7414 14714
rect 7466 14662 7478 14714
rect 7530 14662 7542 14714
rect 7594 14662 7606 14714
rect 7658 14662 10350 14714
rect 10402 14662 10414 14714
rect 10466 14662 10478 14714
rect 10530 14662 10542 14714
rect 10594 14662 10606 14714
rect 10658 14662 13350 14714
rect 13402 14662 13414 14714
rect 13466 14662 13478 14714
rect 13530 14662 13542 14714
rect 13594 14662 13606 14714
rect 13658 14662 16350 14714
rect 16402 14662 16414 14714
rect 16466 14662 16478 14714
rect 16530 14662 16542 14714
rect 16594 14662 16606 14714
rect 16658 14662 19350 14714
rect 19402 14662 19414 14714
rect 19466 14662 19478 14714
rect 19530 14662 19542 14714
rect 19594 14662 19606 14714
rect 19658 14662 22350 14714
rect 22402 14662 22414 14714
rect 22466 14662 22478 14714
rect 22530 14662 22542 14714
rect 22594 14662 22606 14714
rect 22658 14662 24012 14714
rect 1104 14640 24012 14662
rect 7285 14603 7343 14609
rect 1688 14572 7052 14600
rect 1688 14405 1716 14572
rect 2409 14535 2467 14541
rect 2409 14501 2421 14535
rect 2455 14501 2467 14535
rect 3789 14535 3847 14541
rect 2409 14495 2467 14501
rect 2746 14504 3096 14532
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2424 14396 2452 14495
rect 2746 14476 2774 14504
rect 2682 14424 2688 14476
rect 2740 14436 2774 14476
rect 2740 14424 2746 14436
rect 2958 14424 2964 14476
rect 3016 14424 3022 14476
rect 2179 14368 2452 14396
rect 2777 14399 2835 14405
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 2866 14396 2872 14408
rect 2823 14368 2872 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3068 14328 3096 14504
rect 3789 14501 3801 14535
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14396 3663 14399
rect 3804 14396 3832 14495
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4890 14464 4896 14476
rect 4479 14436 4896 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 3651 14368 3832 14396
rect 3651 14365 3663 14368
rect 3605 14359 3663 14365
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4672 14368 5181 14396
rect 4672 14356 4678 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5718 14356 5724 14408
rect 5776 14356 5782 14408
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14396 6239 14399
rect 6546 14396 6552 14408
rect 6227 14368 6552 14396
rect 6227 14365 6239 14368
rect 6181 14359 6239 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 7024 14328 7052 14572
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7374 14600 7380 14612
rect 7331 14572 7380 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 7374 14560 7380 14572
rect 7432 14600 7438 14612
rect 7742 14600 7748 14612
rect 7432 14572 7748 14600
rect 7432 14560 7438 14572
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 9398 14560 9404 14612
rect 9456 14600 9462 14612
rect 9769 14603 9827 14609
rect 9769 14600 9781 14603
rect 9456 14572 9781 14600
rect 9456 14560 9462 14572
rect 9769 14569 9781 14572
rect 9815 14569 9827 14603
rect 9769 14563 9827 14569
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10321 14603 10379 14609
rect 10321 14600 10333 14603
rect 10100 14572 10333 14600
rect 10100 14560 10106 14572
rect 10321 14569 10333 14572
rect 10367 14569 10379 14603
rect 10321 14563 10379 14569
rect 11977 14603 12035 14609
rect 11977 14569 11989 14603
rect 12023 14600 12035 14603
rect 12894 14600 12900 14612
rect 12023 14572 12900 14600
rect 12023 14569 12035 14572
rect 11977 14563 12035 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 13909 14603 13967 14609
rect 13909 14600 13921 14603
rect 13780 14572 13921 14600
rect 13780 14560 13786 14572
rect 13909 14569 13921 14572
rect 13955 14569 13967 14603
rect 13909 14563 13967 14569
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 12434 14532 12440 14544
rect 11848 14504 12440 14532
rect 11848 14492 11854 14504
rect 12434 14492 12440 14504
rect 12492 14492 12498 14544
rect 9122 14424 9128 14476
rect 9180 14424 9186 14476
rect 9217 14467 9275 14473
rect 9217 14433 9229 14467
rect 9263 14464 9275 14467
rect 9582 14464 9588 14476
rect 9263 14436 9588 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 9784 14436 10609 14464
rect 7098 14356 7104 14408
rect 7156 14356 7162 14408
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 8398 14399 8456 14405
rect 8398 14396 8410 14399
rect 7248 14368 8410 14396
rect 7248 14356 7254 14368
rect 8398 14365 8410 14368
rect 8444 14365 8456 14399
rect 8398 14359 8456 14365
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 8754 14396 8760 14408
rect 8711 14368 8760 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 8754 14356 8760 14368
rect 8812 14396 8818 14408
rect 9784 14396 9812 14436
rect 10597 14433 10609 14436
rect 10643 14433 10655 14467
rect 13924 14464 13952 14563
rect 14458 14560 14464 14612
rect 14516 14600 14522 14612
rect 14829 14603 14887 14609
rect 14829 14600 14841 14603
rect 14516 14572 14841 14600
rect 14516 14560 14522 14572
rect 14829 14569 14841 14572
rect 14875 14569 14887 14603
rect 14829 14563 14887 14569
rect 15562 14560 15568 14612
rect 15620 14560 15626 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 18288 14572 18705 14600
rect 18288 14560 18294 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 14550 14492 14556 14544
rect 14608 14532 14614 14544
rect 15013 14535 15071 14541
rect 15013 14532 15025 14535
rect 14608 14504 15025 14532
rect 14608 14492 14614 14504
rect 15013 14501 15025 14504
rect 15059 14501 15071 14535
rect 15013 14495 15071 14501
rect 16942 14492 16948 14544
rect 17000 14532 17006 14544
rect 17000 14504 17356 14532
rect 17000 14492 17006 14504
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 13924 14436 14197 14464
rect 10597 14427 10655 14433
rect 14185 14433 14197 14436
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 8812 14368 9812 14396
rect 9953 14399 10011 14405
rect 8812 14356 8818 14368
rect 9953 14365 9965 14399
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 9214 14328 9220 14340
rect 2884 14300 4200 14328
rect 7024 14300 9220 14328
rect 750 14220 756 14272
rect 808 14260 814 14272
rect 1489 14263 1547 14269
rect 1489 14260 1501 14263
rect 808 14232 1501 14260
rect 808 14220 814 14232
rect 1489 14229 1501 14232
rect 1535 14229 1547 14263
rect 1489 14223 1547 14229
rect 1854 14220 1860 14272
rect 1912 14260 1918 14272
rect 2884 14269 2912 14300
rect 4172 14272 4200 14300
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 9968 14328 9996 14359
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10284 14368 10517 14396
rect 10284 14356 10290 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10612 14396 10640 14427
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 14332 14436 15332 14464
rect 14332 14424 14338 14436
rect 12802 14405 12808 14408
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 10612 14368 12541 14396
rect 10505 14359 10563 14365
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12796 14396 12808 14405
rect 12763 14368 12808 14396
rect 12529 14359 12587 14365
rect 12796 14359 12808 14368
rect 12802 14356 12808 14359
rect 12860 14356 12866 14408
rect 15304 14405 15332 14436
rect 16022 14424 16028 14476
rect 16080 14424 16086 14476
rect 16114 14424 16120 14476
rect 16172 14424 16178 14476
rect 17034 14424 17040 14476
rect 17092 14424 17098 14476
rect 17328 14473 17356 14504
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14433 17371 14467
rect 18708 14464 18736 14563
rect 18874 14560 18880 14612
rect 18932 14600 18938 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 18932 14572 19257 14600
rect 18932 14560 18938 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 19245 14563 19303 14569
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 20990 14560 20996 14612
rect 21048 14560 21054 14612
rect 23106 14560 23112 14612
rect 23164 14600 23170 14612
rect 23293 14603 23351 14609
rect 23293 14600 23305 14603
rect 23164 14572 23305 14600
rect 23164 14560 23170 14572
rect 23293 14569 23305 14572
rect 23339 14569 23351 14603
rect 23293 14563 23351 14569
rect 21910 14532 21916 14544
rect 21652 14504 21916 14532
rect 21652 14473 21680 14504
rect 21910 14492 21916 14504
rect 21968 14492 21974 14544
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 18708 14436 19809 14464
rect 17313 14427 17371 14433
rect 19797 14433 19809 14436
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14433 21695 14467
rect 21637 14427 21695 14433
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14365 15255 14399
rect 15197 14359 15255 14365
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 9692 14300 9996 14328
rect 10864 14331 10922 14337
rect 1949 14263 2007 14269
rect 1949 14260 1961 14263
rect 1912 14232 1961 14260
rect 1912 14220 1918 14232
rect 1949 14229 1961 14232
rect 1995 14229 2007 14263
rect 1949 14223 2007 14229
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14229 2927 14263
rect 2869 14223 2927 14229
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14260 3479 14263
rect 3510 14260 3516 14272
rect 3467 14232 3516 14260
rect 3467 14229 3479 14232
rect 3421 14223 3479 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 4154 14220 4160 14272
rect 4212 14220 4218 14272
rect 4249 14263 4307 14269
rect 4249 14229 4261 14263
rect 4295 14260 4307 14263
rect 4617 14263 4675 14269
rect 4617 14260 4629 14263
rect 4295 14232 4629 14260
rect 4295 14229 4307 14232
rect 4249 14223 4307 14229
rect 4617 14229 4629 14232
rect 4663 14229 4675 14263
rect 4617 14223 4675 14229
rect 5534 14220 5540 14272
rect 5592 14220 5598 14272
rect 5997 14263 6055 14269
rect 5997 14229 6009 14263
rect 6043 14260 6055 14263
rect 6178 14260 6184 14272
rect 6043 14232 6184 14260
rect 6043 14229 6055 14232
rect 5997 14223 6055 14229
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 6549 14263 6607 14269
rect 6549 14229 6561 14263
rect 6595 14260 6607 14263
rect 6914 14260 6920 14272
rect 6595 14232 6920 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 9692 14269 9720 14300
rect 10864 14297 10876 14331
rect 10910 14328 10922 14331
rect 11514 14328 11520 14340
rect 10910 14300 11520 14328
rect 10910 14297 10922 14300
rect 10864 14291 10922 14297
rect 11514 14288 11520 14300
rect 11572 14288 11578 14340
rect 13814 14328 13820 14340
rect 12406 14300 13820 14328
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 7064 14232 9321 14260
rect 7064 14220 7070 14232
rect 9309 14229 9321 14232
rect 9355 14229 9367 14263
rect 9309 14223 9367 14229
rect 9677 14263 9735 14269
rect 9677 14229 9689 14263
rect 9723 14229 9735 14263
rect 9677 14223 9735 14229
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 12406 14260 12434 14300
rect 13814 14288 13820 14300
rect 13872 14328 13878 14340
rect 14642 14328 14648 14340
rect 13872 14300 14648 14328
rect 13872 14288 13878 14300
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 15212 14328 15240 14359
rect 17218 14356 17224 14408
rect 17276 14396 17282 14408
rect 17569 14399 17627 14405
rect 17569 14396 17581 14399
rect 17276 14368 17581 14396
rect 17276 14356 17282 14368
rect 17569 14365 17581 14368
rect 17615 14365 17627 14399
rect 17569 14359 17627 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20806 14396 20812 14408
rect 20211 14368 20812 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21818 14356 21824 14408
rect 21876 14396 21882 14408
rect 21913 14399 21971 14405
rect 21913 14396 21925 14399
rect 21876 14368 21925 14396
rect 21876 14356 21882 14368
rect 21913 14365 21925 14368
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 22462 14356 22468 14408
rect 22520 14396 22526 14408
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 22520 14368 23397 14396
rect 22520 14356 22526 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 15933 14331 15991 14337
rect 15212 14300 15332 14328
rect 15304 14272 15332 14300
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16393 14331 16451 14337
rect 16393 14328 16405 14331
rect 15979 14300 16405 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16393 14297 16405 14300
rect 16439 14297 16451 14331
rect 16393 14291 16451 14297
rect 21450 14288 21456 14340
rect 21508 14328 21514 14340
rect 22158 14331 22216 14337
rect 22158 14328 22170 14331
rect 21508 14300 22170 14328
rect 21508 14288 21514 14300
rect 22158 14297 22170 14300
rect 22204 14297 22216 14331
rect 22158 14291 22216 14297
rect 11112 14232 12434 14260
rect 11112 14220 11118 14232
rect 15286 14220 15292 14272
rect 15344 14220 15350 14272
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14260 15531 14263
rect 15838 14260 15844 14272
rect 15519 14232 15844 14260
rect 15519 14229 15531 14232
rect 15473 14223 15531 14229
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 23566 14220 23572 14272
rect 23624 14220 23630 14272
rect 1104 14170 24164 14192
rect 1104 14118 2850 14170
rect 2902 14118 2914 14170
rect 2966 14118 2978 14170
rect 3030 14118 3042 14170
rect 3094 14118 3106 14170
rect 3158 14118 5850 14170
rect 5902 14118 5914 14170
rect 5966 14118 5978 14170
rect 6030 14118 6042 14170
rect 6094 14118 6106 14170
rect 6158 14118 8850 14170
rect 8902 14118 8914 14170
rect 8966 14118 8978 14170
rect 9030 14118 9042 14170
rect 9094 14118 9106 14170
rect 9158 14118 11850 14170
rect 11902 14118 11914 14170
rect 11966 14118 11978 14170
rect 12030 14118 12042 14170
rect 12094 14118 12106 14170
rect 12158 14118 14850 14170
rect 14902 14118 14914 14170
rect 14966 14118 14978 14170
rect 15030 14118 15042 14170
rect 15094 14118 15106 14170
rect 15158 14118 17850 14170
rect 17902 14118 17914 14170
rect 17966 14118 17978 14170
rect 18030 14118 18042 14170
rect 18094 14118 18106 14170
rect 18158 14118 20850 14170
rect 20902 14118 20914 14170
rect 20966 14118 20978 14170
rect 21030 14118 21042 14170
rect 21094 14118 21106 14170
rect 21158 14118 23850 14170
rect 23902 14118 23914 14170
rect 23966 14118 23978 14170
rect 24030 14118 24042 14170
rect 24094 14118 24106 14170
rect 24158 14118 24164 14170
rect 1104 14096 24164 14118
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 4062 14056 4068 14068
rect 3007 14028 4068 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 4212 14028 5089 14056
rect 4212 14016 4218 14028
rect 5077 14025 5089 14028
rect 5123 14025 5135 14059
rect 5077 14019 5135 14025
rect 6546 14016 6552 14068
rect 6604 14016 6610 14068
rect 6914 14016 6920 14068
rect 6972 14016 6978 14068
rect 7006 14016 7012 14068
rect 7064 14016 7070 14068
rect 8294 14056 8300 14068
rect 7576 14028 8300 14056
rect 2774 13988 2780 14000
rect 1596 13960 2780 13988
rect 1596 13929 1624 13960
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 3418 13948 3424 14000
rect 3476 13988 3482 14000
rect 3476 13960 4752 13988
rect 3476 13948 3482 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 1670 13920 1676 13932
rect 1627 13892 1676 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 1854 13929 1860 13932
rect 1848 13920 1860 13929
rect 1815 13892 1860 13920
rect 1848 13883 1860 13892
rect 1854 13880 1860 13883
rect 1912 13880 1918 13932
rect 2792 13920 2820 13948
rect 3510 13929 3516 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 2792 13892 3249 13920
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3504 13920 3516 13929
rect 3471 13892 3516 13920
rect 3237 13883 3295 13889
rect 3504 13883 3516 13892
rect 3510 13880 3516 13883
rect 3568 13880 3574 13932
rect 4614 13744 4620 13796
rect 4672 13744 4678 13796
rect 4724 13793 4752 13960
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13920 5227 13923
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 5215 13892 5549 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 5537 13889 5549 13892
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 7374 13880 7380 13932
rect 7432 13880 7438 13932
rect 7576 13929 7604 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 9214 14016 9220 14068
rect 9272 14056 9278 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 9272 14028 9321 14056
rect 9272 14016 9278 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 9309 14019 9367 14025
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 9548 14028 10517 14056
rect 9548 14016 9554 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 13780 14028 13829 14056
rect 13780 14016 13786 14028
rect 13817 14025 13829 14028
rect 13863 14025 13875 14059
rect 13817 14019 13875 14025
rect 15194 14016 15200 14068
rect 15252 14016 15258 14068
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 22462 14056 22468 14068
rect 15896 14028 22468 14056
rect 15896 14016 15902 14028
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 22557 14059 22615 14065
rect 22557 14025 22569 14059
rect 22603 14025 22615 14059
rect 22557 14019 22615 14025
rect 12526 13948 12532 14000
rect 12584 13948 12590 14000
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15344 13960 16712 13988
rect 15344 13948 15350 13960
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9263 13892 9505 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 10686 13880 10692 13932
rect 10744 13880 10750 13932
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 13964 13892 14933 13920
rect 13964 13880 13970 13892
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15378 13880 15384 13932
rect 15436 13880 15442 13932
rect 16684 13929 16712 13960
rect 20806 13948 20812 14000
rect 20864 13988 20870 14000
rect 22189 13991 22247 13997
rect 22189 13988 22201 13991
rect 20864 13960 22201 13988
rect 20864 13948 20870 13960
rect 22189 13957 22201 13960
rect 22235 13957 22247 13991
rect 22189 13951 22247 13957
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 21082 13920 21088 13932
rect 20211 13892 21088 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 22572 13920 22600 14019
rect 22922 14016 22928 14068
rect 22980 14056 22986 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22980 14028 23397 14056
rect 22980 14016 22986 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 23569 13923 23627 13929
rect 23569 13920 23581 13923
rect 22572 13892 23581 13920
rect 23569 13889 23581 13892
rect 23615 13889 23627 13923
rect 23569 13883 23627 13889
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5408 13824 6101 13852
rect 5408 13812 5414 13824
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13852 7251 13855
rect 7926 13852 7932 13864
rect 7239 13824 7932 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 8128 13824 8309 13852
rect 4709 13787 4767 13793
rect 4709 13753 4721 13787
rect 4755 13753 4767 13787
rect 4709 13747 4767 13753
rect 4798 13744 4804 13796
rect 4856 13784 4862 13796
rect 7834 13784 7840 13796
rect 4856 13756 7840 13784
rect 4856 13744 4862 13756
rect 7834 13744 7840 13756
rect 7892 13784 7898 13796
rect 8021 13787 8079 13793
rect 8021 13784 8033 13787
rect 7892 13756 8033 13784
rect 7892 13744 7898 13756
rect 8021 13753 8033 13756
rect 8067 13753 8079 13787
rect 8021 13747 8079 13753
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 4632 13716 4660 13744
rect 4212 13688 4660 13716
rect 4212 13676 4218 13688
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 6638 13716 6644 13728
rect 5316 13688 6644 13716
rect 5316 13676 5322 13688
rect 6638 13676 6644 13688
rect 6696 13676 6702 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 8128 13716 8156 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8386 13812 8392 13864
rect 8444 13861 8450 13864
rect 8444 13855 8472 13861
rect 8460 13821 8472 13855
rect 8444 13815 8472 13821
rect 8444 13812 8450 13815
rect 8570 13812 8576 13864
rect 8628 13812 8634 13864
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20772 13824 20821 13852
rect 20772 13812 20778 13824
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 21361 13855 21419 13861
rect 21361 13852 21373 13855
rect 21324 13824 21373 13852
rect 21324 13812 21330 13824
rect 21361 13821 21373 13824
rect 21407 13852 21419 13855
rect 21910 13852 21916 13864
rect 21407 13824 21916 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 21910 13812 21916 13824
rect 21968 13812 21974 13864
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 22097 13855 22155 13861
rect 22097 13821 22109 13855
rect 22143 13852 22155 13855
rect 22649 13855 22707 13861
rect 22649 13852 22661 13855
rect 22143 13824 22661 13852
rect 22143 13821 22155 13824
rect 22097 13815 22155 13821
rect 22649 13821 22661 13824
rect 22695 13821 22707 13855
rect 22649 13815 22707 13821
rect 16853 13787 16911 13793
rect 16853 13753 16865 13787
rect 16899 13784 16911 13787
rect 17770 13784 17776 13796
rect 16899 13756 17776 13784
rect 16899 13753 16911 13756
rect 16853 13747 16911 13753
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 22020 13784 22048 13815
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 23201 13855 23259 13861
rect 23201 13852 23213 13855
rect 23072 13824 23213 13852
rect 23072 13812 23078 13824
rect 23201 13821 23213 13824
rect 23247 13821 23259 13855
rect 23201 13815 23259 13821
rect 22020 13756 22094 13784
rect 22066 13728 22094 13756
rect 7156 13688 8156 13716
rect 7156 13676 7162 13688
rect 14366 13676 14372 13728
rect 14424 13676 14430 13728
rect 20717 13719 20775 13725
rect 20717 13685 20729 13719
rect 20763 13716 20775 13719
rect 21358 13716 21364 13728
rect 20763 13688 21364 13716
rect 20763 13685 20775 13688
rect 20717 13679 20775 13685
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 22066 13688 22100 13728
rect 22094 13676 22100 13688
rect 22152 13716 22158 13728
rect 22830 13716 22836 13728
rect 22152 13688 22836 13716
rect 22152 13676 22158 13688
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 1104 13626 24012 13648
rect 1104 13574 1350 13626
rect 1402 13574 1414 13626
rect 1466 13574 1478 13626
rect 1530 13574 1542 13626
rect 1594 13574 1606 13626
rect 1658 13574 4350 13626
rect 4402 13574 4414 13626
rect 4466 13574 4478 13626
rect 4530 13574 4542 13626
rect 4594 13574 4606 13626
rect 4658 13574 7350 13626
rect 7402 13574 7414 13626
rect 7466 13574 7478 13626
rect 7530 13574 7542 13626
rect 7594 13574 7606 13626
rect 7658 13574 10350 13626
rect 10402 13574 10414 13626
rect 10466 13574 10478 13626
rect 10530 13574 10542 13626
rect 10594 13574 10606 13626
rect 10658 13574 13350 13626
rect 13402 13574 13414 13626
rect 13466 13574 13478 13626
rect 13530 13574 13542 13626
rect 13594 13574 13606 13626
rect 13658 13574 16350 13626
rect 16402 13574 16414 13626
rect 16466 13574 16478 13626
rect 16530 13574 16542 13626
rect 16594 13574 16606 13626
rect 16658 13574 19350 13626
rect 19402 13574 19414 13626
rect 19466 13574 19478 13626
rect 19530 13574 19542 13626
rect 19594 13574 19606 13626
rect 19658 13574 22350 13626
rect 22402 13574 22414 13626
rect 22466 13574 22478 13626
rect 22530 13574 22542 13626
rect 22594 13574 22606 13626
rect 22658 13574 24012 13626
rect 1104 13552 24012 13574
rect 1670 13512 1676 13524
rect 1504 13484 1676 13512
rect 1504 13385 1532 13484
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4706 13512 4712 13524
rect 4304 13484 4712 13512
rect 4304 13472 4310 13484
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 5629 13515 5687 13521
rect 5629 13481 5641 13515
rect 5675 13512 5687 13515
rect 5718 13512 5724 13524
rect 5675 13484 5724 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 7156 13484 7297 13512
rect 7156 13472 7162 13484
rect 7285 13481 7297 13484
rect 7331 13481 7343 13515
rect 7285 13475 7343 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12492 13484 12633 13512
rect 12492 13472 12498 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 13262 13512 13268 13524
rect 13136 13484 13268 13512
rect 13136 13472 13142 13484
rect 13262 13472 13268 13484
rect 13320 13512 13326 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13320 13484 13645 13512
rect 13320 13472 13326 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 20806 13472 20812 13524
rect 20864 13472 20870 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 23293 13515 23351 13521
rect 23293 13512 23305 13515
rect 21140 13484 23305 13512
rect 21140 13472 21146 13484
rect 23293 13481 23305 13484
rect 23339 13512 23351 13515
rect 23474 13512 23480 13524
rect 23339 13484 23480 13512
rect 23339 13481 23351 13484
rect 23293 13475 23351 13481
rect 23474 13472 23480 13484
rect 23532 13472 23538 13524
rect 2869 13447 2927 13453
rect 2869 13413 2881 13447
rect 2915 13444 2927 13447
rect 11057 13447 11115 13453
rect 2915 13416 4568 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 3620 13385 3648 13416
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13345 1547 13379
rect 1489 13339 1547 13345
rect 3605 13379 3663 13385
rect 3605 13345 3617 13379
rect 3651 13345 3663 13379
rect 3605 13339 3663 13345
rect 3789 13379 3847 13385
rect 3789 13345 3801 13379
rect 3835 13376 3847 13379
rect 4154 13376 4160 13388
rect 3835 13348 4160 13376
rect 3835 13345 3847 13348
rect 3789 13339 3847 13345
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 4396 13348 4445 13376
rect 4396 13336 4402 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 4540 13376 4568 13416
rect 11057 13413 11069 13447
rect 11103 13444 11115 13447
rect 13170 13444 13176 13456
rect 11103 13416 13176 13444
rect 11103 13413 11115 13416
rect 11057 13407 11115 13413
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 15381 13447 15439 13453
rect 15381 13413 15393 13447
rect 15427 13413 15439 13447
rect 15381 13407 15439 13413
rect 4826 13379 4884 13385
rect 4826 13376 4838 13379
rect 4540 13348 4838 13376
rect 4433 13339 4491 13345
rect 4826 13345 4838 13348
rect 4872 13345 4884 13379
rect 4826 13339 4884 13345
rect 4982 13336 4988 13388
rect 5040 13376 5046 13388
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 5040 13348 6040 13376
rect 5040 13336 5046 13348
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3936 13280 3985 13308
rect 3936 13268 3942 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 1756 13243 1814 13249
rect 1756 13209 1768 13243
rect 1802 13240 1814 13243
rect 1854 13240 1860 13252
rect 1802 13212 1860 13240
rect 1802 13209 1814 13212
rect 1756 13203 1814 13209
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 2590 13200 2596 13252
rect 2648 13240 2654 13252
rect 2961 13243 3019 13249
rect 2961 13240 2973 13243
rect 2648 13212 2973 13240
rect 2648 13200 2654 13212
rect 2961 13209 2973 13212
rect 3007 13209 3019 13243
rect 2961 13203 3019 13209
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 5920 13172 5948 13271
rect 6012 13240 6040 13348
rect 6932 13348 7941 13376
rect 6178 13317 6184 13320
rect 6172 13308 6184 13317
rect 6139 13280 6184 13308
rect 6172 13271 6184 13280
rect 6178 13268 6184 13271
rect 6236 13268 6242 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 6932 13308 6960 13348
rect 7929 13345 7941 13348
rect 7975 13376 7987 13379
rect 8110 13376 8116 13388
rect 7975 13348 8116 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 13265 13379 13323 13385
rect 13265 13345 13277 13379
rect 13311 13376 13323 13379
rect 13722 13376 13728 13388
rect 13311 13348 13728 13376
rect 13311 13345 13323 13348
rect 13265 13339 13323 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 6696 13280 6960 13308
rect 6696 13268 6702 13280
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7064 13280 7757 13308
rect 7064 13268 7070 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 8662 13308 8668 13320
rect 7892 13280 8668 13308
rect 7892 13268 7898 13280
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 11146 13268 11152 13320
rect 11204 13268 11210 13320
rect 12342 13268 12348 13320
rect 12400 13268 12406 13320
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 14366 13308 14372 13320
rect 13127 13280 14372 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15396 13308 15424 13407
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 21634 13444 21640 13456
rect 16264 13416 21640 13444
rect 16264 13404 16270 13416
rect 16025 13379 16083 13385
rect 16025 13345 16037 13379
rect 16071 13376 16083 13379
rect 16114 13376 16120 13388
rect 16071 13348 16120 13376
rect 16071 13345 16083 13348
rect 16025 13339 16083 13345
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 18414 13376 18420 13388
rect 17328 13348 18420 13376
rect 15151 13280 15424 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15930 13268 15936 13320
rect 15988 13308 15994 13320
rect 17328 13317 17356 13348
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 20456 13385 20484 13416
rect 21634 13404 21640 13416
rect 21692 13404 21698 13456
rect 20441 13379 20499 13385
rect 20441 13345 20453 13379
rect 20487 13345 20499 13379
rect 20441 13339 20499 13345
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21177 13379 21235 13385
rect 21177 13376 21189 13379
rect 20680 13348 21189 13376
rect 20680 13336 20686 13348
rect 21177 13345 21189 13348
rect 21223 13345 21235 13379
rect 21177 13339 21235 13345
rect 21358 13336 21364 13388
rect 21416 13336 21422 13388
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 15988 13280 16773 13308
rect 15988 13268 15994 13280
rect 16761 13277 16773 13280
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 8570 13240 8576 13252
rect 6012 13212 8576 13240
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 13170 13200 13176 13252
rect 13228 13240 13234 13252
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 13228 13212 13553 13240
rect 13228 13200 13234 13212
rect 13541 13209 13553 13212
rect 13587 13240 13599 13243
rect 15286 13240 15292 13252
rect 13587 13212 15292 13240
rect 13587 13209 13599 13212
rect 13541 13203 13599 13209
rect 15286 13200 15292 13212
rect 15344 13200 15350 13252
rect 15749 13243 15807 13249
rect 15749 13209 15761 13243
rect 15795 13240 15807 13243
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15795 13212 16221 13240
rect 15795 13209 15807 13212
rect 15749 13203 15807 13209
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16776 13240 16804 13271
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17552 13280 17601 13308
rect 17552 13268 17558 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 20530 13308 20536 13320
rect 19751 13280 20536 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21542 13308 21548 13320
rect 21039 13280 21548 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 21818 13268 21824 13320
rect 21876 13308 21882 13320
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21876 13280 21925 13308
rect 21876 13268 21882 13280
rect 21913 13277 21925 13280
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 23382 13268 23388 13320
rect 23440 13268 23446 13320
rect 16776 13212 17632 13240
rect 16209 13203 16267 13209
rect 17604 13184 17632 13212
rect 18782 13200 18788 13252
rect 18840 13240 18846 13252
rect 21174 13240 21180 13252
rect 18840 13212 21180 13240
rect 18840 13200 18846 13212
rect 21174 13200 21180 13212
rect 21232 13200 21238 13252
rect 21453 13243 21511 13249
rect 21453 13209 21465 13243
rect 21499 13240 21511 13243
rect 21634 13240 21640 13252
rect 21499 13212 21640 13240
rect 21499 13209 21511 13212
rect 21453 13203 21511 13209
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22186 13249 22192 13252
rect 22180 13203 22192 13249
rect 22186 13200 22192 13203
rect 22244 13200 22250 13252
rect 4028 13144 5948 13172
rect 4028 13132 4034 13144
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 7834 13132 7840 13184
rect 7892 13132 7898 13184
rect 11330 13132 11336 13184
rect 11388 13132 11394 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 11793 13175 11851 13181
rect 11793 13172 11805 13175
rect 11756 13144 11805 13172
rect 11756 13132 11762 13144
rect 11793 13141 11805 13144
rect 11839 13141 11851 13175
rect 11793 13135 11851 13141
rect 14734 13132 14740 13184
rect 14792 13172 14798 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14792 13144 14933 13172
rect 14792 13132 14798 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 14921 13135 14979 13141
rect 15838 13132 15844 13184
rect 15896 13132 15902 13184
rect 17126 13132 17132 13184
rect 17184 13132 17190 13184
rect 17402 13132 17408 13184
rect 17460 13132 17466 13184
rect 17586 13132 17592 13184
rect 17644 13132 17650 13184
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19521 13175 19579 13181
rect 19521 13172 19533 13175
rect 19484 13144 19533 13172
rect 19484 13132 19490 13144
rect 19521 13141 19533 13144
rect 19567 13141 19579 13175
rect 19521 13135 19579 13141
rect 19886 13132 19892 13184
rect 19944 13132 19950 13184
rect 20254 13132 20260 13184
rect 20312 13132 20318 13184
rect 20349 13175 20407 13181
rect 20349 13141 20361 13175
rect 20395 13172 20407 13175
rect 20622 13172 20628 13184
rect 20395 13144 20628 13172
rect 20395 13141 20407 13144
rect 20349 13135 20407 13141
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 21542 13132 21548 13184
rect 21600 13172 21606 13184
rect 21821 13175 21879 13181
rect 21821 13172 21833 13175
rect 21600 13144 21833 13172
rect 21600 13132 21606 13144
rect 21821 13141 21833 13144
rect 21867 13141 21879 13175
rect 21821 13135 21879 13141
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 22738 13172 22744 13184
rect 21968 13144 22744 13172
rect 21968 13132 21974 13144
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 23569 13175 23627 13181
rect 23569 13141 23581 13175
rect 23615 13172 23627 13175
rect 24302 13172 24308 13184
rect 23615 13144 24308 13172
rect 23615 13141 23627 13144
rect 23569 13135 23627 13141
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 1104 13082 24164 13104
rect 1104 13030 2850 13082
rect 2902 13030 2914 13082
rect 2966 13030 2978 13082
rect 3030 13030 3042 13082
rect 3094 13030 3106 13082
rect 3158 13030 5850 13082
rect 5902 13030 5914 13082
rect 5966 13030 5978 13082
rect 6030 13030 6042 13082
rect 6094 13030 6106 13082
rect 6158 13030 8850 13082
rect 8902 13030 8914 13082
rect 8966 13030 8978 13082
rect 9030 13030 9042 13082
rect 9094 13030 9106 13082
rect 9158 13030 11850 13082
rect 11902 13030 11914 13082
rect 11966 13030 11978 13082
rect 12030 13030 12042 13082
rect 12094 13030 12106 13082
rect 12158 13030 14850 13082
rect 14902 13030 14914 13082
rect 14966 13030 14978 13082
rect 15030 13030 15042 13082
rect 15094 13030 15106 13082
rect 15158 13030 17850 13082
rect 17902 13030 17914 13082
rect 17966 13030 17978 13082
rect 18030 13030 18042 13082
rect 18094 13030 18106 13082
rect 18158 13030 20850 13082
rect 20902 13030 20914 13082
rect 20966 13030 20978 13082
rect 21030 13030 21042 13082
rect 21094 13030 21106 13082
rect 21158 13030 23850 13082
rect 23902 13030 23914 13082
rect 23966 13030 23978 13082
rect 24030 13030 24042 13082
rect 24094 13030 24106 13082
rect 24158 13030 24164 13082
rect 1104 13008 24164 13030
rect 1302 12928 1308 12980
rect 1360 12968 1366 12980
rect 1489 12971 1547 12977
rect 1489 12968 1501 12971
rect 1360 12940 1501 12968
rect 1360 12928 1366 12940
rect 1489 12937 1501 12940
rect 1535 12937 1547 12971
rect 1489 12931 1547 12937
rect 1854 12928 1860 12980
rect 1912 12928 1918 12980
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12937 2191 12971
rect 2133 12931 2191 12937
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2041 12835 2099 12841
rect 1719 12804 1992 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 1964 12628 1992 12804
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2148 12832 2176 12931
rect 2590 12928 2596 12980
rect 2648 12928 2654 12980
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 5350 12968 5356 12980
rect 3936 12940 5356 12968
rect 3936 12928 3942 12940
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 7374 12968 7380 12980
rect 6012 12940 7380 12968
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 2682 12900 2688 12912
rect 2547 12872 2688 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3053 12903 3111 12909
rect 3053 12900 3065 12903
rect 2832 12872 3065 12900
rect 2832 12860 2838 12872
rect 3053 12869 3065 12872
rect 3099 12900 3111 12903
rect 3099 12872 4016 12900
rect 3099 12869 3111 12872
rect 3053 12863 3111 12869
rect 3988 12844 4016 12872
rect 4080 12872 5948 12900
rect 2087 12804 2176 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 3878 12792 3884 12844
rect 3936 12792 3942 12844
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 4080 12764 4108 12872
rect 4240 12835 4298 12841
rect 4240 12801 4252 12835
rect 4286 12832 4298 12835
rect 4522 12832 4528 12844
rect 4286 12804 4528 12832
rect 4286 12801 4298 12804
rect 4240 12795 4298 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 2731 12736 4108 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 5534 12628 5540 12640
rect 1964 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 5920 12628 5948 12872
rect 6012 12841 6040 12940
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 7834 12928 7840 12980
rect 7892 12928 7898 12980
rect 9861 12971 9919 12977
rect 9861 12937 9873 12971
rect 9907 12937 9919 12971
rect 11422 12968 11428 12980
rect 9861 12931 9919 12937
rect 10796 12940 11428 12968
rect 8754 12900 8760 12912
rect 6380 12872 8760 12900
rect 6380 12841 6408 12872
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6621 12835 6679 12841
rect 6621 12832 6633 12835
rect 6365 12795 6423 12801
rect 6472 12804 6633 12832
rect 6472 12764 6500 12804
rect 6621 12801 6633 12804
rect 6667 12801 6679 12835
rect 6621 12795 6679 12801
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9876 12832 9904 12931
rect 9723 12804 9904 12832
rect 10229 12835 10287 12841
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10275 12804 10701 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 6196 12736 6500 12764
rect 6196 12705 6224 12736
rect 6181 12699 6239 12705
rect 6181 12665 6193 12699
rect 6227 12665 6239 12699
rect 6181 12659 6239 12665
rect 7745 12699 7803 12705
rect 7745 12665 7757 12699
rect 7791 12696 7803 12699
rect 8404 12696 8432 12792
rect 7791 12668 8432 12696
rect 7791 12665 7803 12668
rect 7745 12659 7803 12665
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 8720 12668 8769 12696
rect 8720 12656 8726 12668
rect 8757 12665 8769 12668
rect 8803 12665 8815 12699
rect 8956 12696 8984 12795
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10192 12736 10333 12764
rect 10192 12724 10198 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12764 10563 12767
rect 10796 12764 10824 12940
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 12342 12968 12348 12980
rect 11563 12940 12348 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 12989 12971 13047 12977
rect 12989 12968 13001 12971
rect 12860 12940 13001 12968
rect 12860 12928 12866 12940
rect 12989 12937 13001 12940
rect 13035 12937 13047 12971
rect 12989 12931 13047 12937
rect 14292 12940 15792 12968
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 12630 12903 12688 12909
rect 12630 12900 12642 12903
rect 11388 12872 12642 12900
rect 11388 12860 11394 12872
rect 12630 12869 12642 12872
rect 12676 12869 12688 12903
rect 12630 12863 12688 12869
rect 11422 12792 11428 12844
rect 11480 12832 11486 12844
rect 14292 12841 14320 12940
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 15764 12900 15792 12940
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 16715 12940 18644 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16022 12900 16028 12912
rect 14792 12872 14872 12900
rect 15764 12872 16028 12900
rect 14792 12860 14798 12872
rect 14844 12841 14872 12872
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 11480 12804 13185 12832
rect 11480 12792 11486 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14820 12835 14878 12841
rect 14820 12801 14832 12835
rect 14866 12801 14878 12835
rect 14820 12795 14878 12801
rect 17586 12792 17592 12844
rect 17644 12792 17650 12844
rect 18616 12841 18644 12940
rect 18782 12928 18788 12980
rect 18840 12928 18846 12980
rect 19886 12968 19892 12980
rect 19076 12940 19892 12968
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12832 18935 12835
rect 19076 12832 19104 12940
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 20625 12971 20683 12977
rect 20625 12968 20637 12971
rect 20588 12940 20637 12968
rect 20588 12928 20594 12940
rect 20625 12937 20637 12940
rect 20671 12937 20683 12971
rect 20625 12931 20683 12937
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 20993 12971 21051 12977
rect 20993 12968 21005 12971
rect 20772 12940 21005 12968
rect 20772 12928 20778 12940
rect 20993 12937 21005 12940
rect 21039 12937 21051 12971
rect 20993 12931 21051 12937
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 23198 12968 23204 12980
rect 21232 12940 23204 12968
rect 21232 12928 21238 12940
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 21818 12900 21824 12912
rect 19208 12872 21824 12900
rect 19208 12860 19214 12872
rect 21818 12860 21824 12872
rect 21876 12860 21882 12912
rect 19426 12841 19432 12844
rect 19420 12832 19432 12841
rect 18923 12804 19104 12832
rect 19387 12804 19432 12832
rect 18923 12801 18935 12804
rect 18877 12795 18935 12801
rect 19420 12795 19432 12804
rect 19426 12792 19432 12795
rect 19484 12792 19490 12844
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 22462 12792 22468 12844
rect 22520 12792 22526 12844
rect 22738 12792 22744 12844
rect 22796 12792 22802 12844
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 23661 12835 23719 12841
rect 23661 12832 23673 12835
rect 23348 12804 23673 12832
rect 23348 12792 23354 12804
rect 23661 12801 23673 12804
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 10551 12736 10824 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11112 12736 11253 12764
rect 11112 12724 11118 12736
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 12894 12724 12900 12776
rect 12952 12764 12958 12776
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 12952 12736 14565 12764
rect 12952 12724 12958 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 17310 12724 17316 12776
rect 17368 12724 17374 12776
rect 17472 12767 17530 12773
rect 17472 12733 17484 12767
rect 17518 12764 17530 12767
rect 17770 12764 17776 12776
rect 17518 12736 17776 12764
rect 17518 12733 17530 12736
rect 17472 12727 17530 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 17862 12724 17868 12776
rect 17920 12724 17926 12776
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 11790 12696 11796 12708
rect 8956 12668 11796 12696
rect 8757 12659 8815 12665
rect 11790 12656 11796 12668
rect 11848 12656 11854 12708
rect 18230 12656 18236 12708
rect 18288 12696 18294 12708
rect 18524 12696 18552 12727
rect 19150 12724 19156 12776
rect 19208 12724 19214 12776
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 21082 12764 21088 12776
rect 20312 12736 21088 12764
rect 20312 12724 20318 12736
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 21266 12724 21272 12776
rect 21324 12724 21330 12776
rect 22603 12767 22661 12773
rect 22603 12764 22615 12767
rect 21560 12736 22615 12764
rect 18288 12668 18552 12696
rect 20533 12699 20591 12705
rect 18288 12656 18294 12668
rect 20533 12665 20545 12699
rect 20579 12696 20591 12699
rect 21174 12696 21180 12708
rect 20579 12668 21180 12696
rect 20579 12665 20591 12668
rect 20533 12659 20591 12665
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 6638 12628 6644 12640
rect 5920 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9456 12600 9505 12628
rect 9456 12588 9462 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 11514 12588 11520 12640
rect 11572 12628 11578 12640
rect 12986 12628 12992 12640
rect 11572 12600 12992 12628
rect 11572 12588 11578 12600
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 14458 12588 14464 12640
rect 14516 12588 14522 12640
rect 19061 12631 19119 12637
rect 19061 12597 19073 12631
rect 19107 12628 19119 12631
rect 19794 12628 19800 12640
rect 19107 12600 19800 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 21560 12628 21588 12736
rect 22603 12733 22615 12736
rect 22649 12733 22661 12767
rect 22603 12727 22661 12733
rect 22922 12724 22928 12776
rect 22980 12764 22986 12776
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22980 12736 23029 12764
rect 22980 12724 22986 12736
rect 23017 12733 23029 12736
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 23474 12724 23480 12776
rect 23532 12724 23538 12776
rect 21637 12699 21695 12705
rect 21637 12665 21649 12699
rect 21683 12696 21695 12699
rect 21683 12668 22094 12696
rect 21683 12665 21695 12668
rect 21637 12659 21695 12665
rect 22066 12640 22094 12668
rect 21416 12600 21588 12628
rect 21821 12631 21879 12637
rect 21416 12588 21422 12600
rect 21821 12597 21833 12631
rect 21867 12628 21879 12631
rect 21910 12628 21916 12640
rect 21867 12600 21916 12628
rect 21867 12597 21879 12600
rect 21821 12591 21879 12597
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 22066 12600 22100 12640
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 1104 12538 24012 12560
rect 1104 12486 1350 12538
rect 1402 12486 1414 12538
rect 1466 12486 1478 12538
rect 1530 12486 1542 12538
rect 1594 12486 1606 12538
rect 1658 12486 4350 12538
rect 4402 12486 4414 12538
rect 4466 12486 4478 12538
rect 4530 12486 4542 12538
rect 4594 12486 4606 12538
rect 4658 12486 7350 12538
rect 7402 12486 7414 12538
rect 7466 12486 7478 12538
rect 7530 12486 7542 12538
rect 7594 12486 7606 12538
rect 7658 12486 10350 12538
rect 10402 12486 10414 12538
rect 10466 12486 10478 12538
rect 10530 12486 10542 12538
rect 10594 12486 10606 12538
rect 10658 12486 13350 12538
rect 13402 12486 13414 12538
rect 13466 12486 13478 12538
rect 13530 12486 13542 12538
rect 13594 12486 13606 12538
rect 13658 12486 16350 12538
rect 16402 12486 16414 12538
rect 16466 12486 16478 12538
rect 16530 12486 16542 12538
rect 16594 12486 16606 12538
rect 16658 12486 19350 12538
rect 19402 12486 19414 12538
rect 19466 12486 19478 12538
rect 19530 12486 19542 12538
rect 19594 12486 19606 12538
rect 19658 12486 22350 12538
rect 22402 12486 22414 12538
rect 22466 12486 22478 12538
rect 22530 12486 22542 12538
rect 22594 12486 22606 12538
rect 22658 12486 24012 12538
rect 1104 12464 24012 12486
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12424 3663 12427
rect 4246 12424 4252 12436
rect 3651 12396 4252 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 10134 12424 10140 12436
rect 9140 12396 10140 12424
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12356 1639 12359
rect 9140 12356 9168 12396
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 11422 12424 11428 12436
rect 10643 12396 11428 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 14369 12427 14427 12433
rect 11572 12396 11744 12424
rect 11572 12384 11578 12396
rect 1627 12328 9168 12356
rect 10505 12359 10563 12365
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 10505 12325 10517 12359
rect 10551 12325 10563 12359
rect 11716 12356 11744 12396
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 14415 12396 15792 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 11790 12356 11796 12368
rect 11716 12328 11796 12356
rect 10505 12319 10563 12325
rect 10520 12288 10548 12319
rect 11790 12316 11796 12328
rect 11848 12356 11854 12368
rect 11848 12328 12848 12356
rect 11848 12316 11854 12328
rect 11054 12288 11060 12300
rect 10520 12260 11060 12288
rect 11054 12248 11060 12260
rect 11112 12288 11118 12300
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11112 12260 11529 12288
rect 11112 12248 11118 12260
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12342 12288 12348 12300
rect 12299 12260 12348 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 382 12180 388 12232
rect 440 12220 446 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 440 12192 1409 12220
rect 440 12180 446 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 3418 12180 3424 12232
rect 3476 12180 3482 12232
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8662 12220 8668 12232
rect 8619 12192 8668 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8812 12192 9137 12220
rect 8812 12180 8818 12192
rect 9125 12189 9137 12192
rect 9171 12220 9183 12223
rect 9214 12220 9220 12232
rect 9171 12192 9220 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 9398 12229 9404 12232
rect 9392 12183 9404 12229
rect 9398 12180 9404 12183
rect 9456 12180 9462 12232
rect 11238 12180 11244 12232
rect 11296 12180 11302 12232
rect 11422 12229 11428 12232
rect 11400 12223 11428 12229
rect 11400 12189 11412 12223
rect 11400 12183 11428 12189
rect 11422 12180 11428 12183
rect 11480 12180 11486 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 12483 12192 12572 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 12544 12096 12572 12192
rect 12820 12152 12848 12328
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 13924 12260 14565 12288
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13924 12229 13952 12260
rect 14553 12257 14565 12260
rect 14599 12257 14611 12291
rect 15764 12288 15792 12396
rect 16022 12384 16028 12436
rect 16080 12384 16086 12436
rect 16574 12424 16580 12436
rect 16500 12396 16580 12424
rect 15933 12359 15991 12365
rect 15933 12325 15945 12359
rect 15979 12356 15991 12359
rect 16500 12356 16528 12396
rect 16574 12384 16580 12396
rect 16632 12424 16638 12436
rect 17770 12424 17776 12436
rect 16632 12396 17776 12424
rect 16632 12384 16638 12396
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 18325 12427 18383 12433
rect 18325 12393 18337 12427
rect 18371 12424 18383 12427
rect 18414 12424 18420 12436
rect 18371 12396 18420 12424
rect 18371 12393 18383 12396
rect 18325 12387 18383 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 20714 12384 20720 12436
rect 20772 12384 20778 12436
rect 21729 12427 21787 12433
rect 21729 12393 21741 12427
rect 21775 12424 21787 12427
rect 22186 12424 22192 12436
rect 21775 12396 22192 12424
rect 21775 12393 21787 12396
rect 21729 12387 21787 12393
rect 22186 12384 22192 12396
rect 22244 12384 22250 12436
rect 23201 12427 23259 12433
rect 23201 12393 23213 12427
rect 23247 12424 23259 12427
rect 23290 12424 23296 12436
rect 23247 12396 23296 12424
rect 23247 12393 23259 12396
rect 23201 12387 23259 12393
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 15979 12328 16528 12356
rect 20625 12359 20683 12365
rect 15979 12325 15991 12328
rect 15933 12319 15991 12325
rect 20625 12325 20637 12359
rect 20671 12325 20683 12359
rect 20625 12319 20683 12325
rect 16206 12288 16212 12300
rect 15764 12260 16212 12288
rect 14553 12251 14611 12257
rect 16206 12248 16212 12260
rect 16264 12288 16270 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16264 12260 16589 12288
rect 16264 12248 16270 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 18969 12291 19027 12297
rect 18969 12257 18981 12291
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 13909 12223 13967 12229
rect 13909 12220 13921 12223
rect 12952 12192 13921 12220
rect 12952 12180 12958 12192
rect 13909 12189 13921 12192
rect 13955 12189 13967 12223
rect 13909 12183 13967 12189
rect 14090 12180 14096 12232
rect 14148 12220 14154 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 14148 12192 14197 12220
rect 14148 12180 14154 12192
rect 14185 12189 14197 12192
rect 14231 12189 14243 12223
rect 14185 12183 14243 12189
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 14809 12223 14867 12229
rect 14809 12220 14821 12223
rect 14516 12192 14821 12220
rect 14516 12180 14522 12192
rect 14809 12189 14821 12192
rect 14855 12189 14867 12223
rect 14809 12183 14867 12189
rect 16850 12180 16856 12232
rect 16908 12180 16914 12232
rect 17126 12229 17132 12232
rect 17120 12183 17132 12229
rect 17126 12180 17132 12183
rect 17184 12180 17190 12232
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 18984 12220 19012 12251
rect 19150 12248 19156 12300
rect 19208 12288 19214 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19208 12260 19257 12288
rect 19208 12248 19214 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 20640 12288 20668 12319
rect 23566 12316 23572 12368
rect 23624 12316 23630 12368
rect 21358 12288 21364 12300
rect 20640 12260 21364 12288
rect 19245 12251 19303 12257
rect 21358 12248 21364 12260
rect 21416 12248 21422 12300
rect 21818 12248 21824 12300
rect 21876 12248 21882 12300
rect 17736 12192 19012 12220
rect 17736 12180 17742 12192
rect 12820 12124 13124 12152
rect 13096 12096 13124 12124
rect 13262 12112 13268 12164
rect 13320 12152 13326 12164
rect 13642 12155 13700 12161
rect 13642 12152 13654 12155
rect 13320 12124 13654 12152
rect 13320 12112 13326 12124
rect 13642 12121 13654 12124
rect 13688 12121 13700 12155
rect 13642 12115 13700 12121
rect 15838 12112 15844 12164
rect 15896 12152 15902 12164
rect 16393 12155 16451 12161
rect 16393 12152 16405 12155
rect 15896 12124 16405 12152
rect 15896 12112 15902 12124
rect 16393 12121 16405 12124
rect 16439 12152 16451 12155
rect 18984 12152 19012 12192
rect 19512 12223 19570 12229
rect 19512 12189 19524 12223
rect 19558 12220 19570 12223
rect 19794 12220 19800 12232
rect 19558 12192 19800 12220
rect 19558 12189 19570 12192
rect 19512 12183 19570 12189
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 21542 12180 21548 12232
rect 21600 12180 21606 12232
rect 22094 12229 22100 12232
rect 22088 12220 22100 12229
rect 22055 12192 22100 12220
rect 22088 12183 22100 12192
rect 22094 12180 22100 12183
rect 22152 12180 22158 12232
rect 23198 12180 23204 12232
rect 23256 12220 23262 12232
rect 23385 12223 23443 12229
rect 23385 12220 23397 12223
rect 23256 12192 23397 12220
rect 23256 12180 23262 12192
rect 23385 12189 23397 12192
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 22830 12152 22836 12164
rect 16439 12124 18736 12152
rect 18984 12124 22836 12152
rect 16439 12121 16451 12124
rect 16393 12115 16451 12121
rect 18708 12096 18736 12124
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12084 8815 12087
rect 9398 12084 9404 12096
rect 8803 12056 9404 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 12526 12044 12532 12096
rect 12584 12044 12590 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 15286 12084 15292 12096
rect 13136 12056 15292 12084
rect 13136 12044 13142 12056
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 16482 12044 16488 12096
rect 16540 12044 16546 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18598 12084 18604 12096
rect 18288 12056 18604 12084
rect 18288 12044 18294 12056
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 18690 12044 18696 12096
rect 18748 12044 18754 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 19242 12084 19248 12096
rect 18831 12056 19248 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 21082 12044 21088 12096
rect 21140 12084 21146 12096
rect 21634 12084 21640 12096
rect 21140 12056 21640 12084
rect 21140 12044 21146 12056
rect 21634 12044 21640 12056
rect 21692 12084 21698 12096
rect 22186 12084 22192 12096
rect 21692 12056 22192 12084
rect 21692 12044 21698 12056
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 1104 11994 24164 12016
rect 1104 11942 2850 11994
rect 2902 11942 2914 11994
rect 2966 11942 2978 11994
rect 3030 11942 3042 11994
rect 3094 11942 3106 11994
rect 3158 11942 5850 11994
rect 5902 11942 5914 11994
rect 5966 11942 5978 11994
rect 6030 11942 6042 11994
rect 6094 11942 6106 11994
rect 6158 11942 8850 11994
rect 8902 11942 8914 11994
rect 8966 11942 8978 11994
rect 9030 11942 9042 11994
rect 9094 11942 9106 11994
rect 9158 11942 11850 11994
rect 11902 11942 11914 11994
rect 11966 11942 11978 11994
rect 12030 11942 12042 11994
rect 12094 11942 12106 11994
rect 12158 11942 14850 11994
rect 14902 11942 14914 11994
rect 14966 11942 14978 11994
rect 15030 11942 15042 11994
rect 15094 11942 15106 11994
rect 15158 11942 17850 11994
rect 17902 11942 17914 11994
rect 17966 11942 17978 11994
rect 18030 11942 18042 11994
rect 18094 11942 18106 11994
rect 18158 11942 20850 11994
rect 20902 11942 20914 11994
rect 20966 11942 20978 11994
rect 21030 11942 21042 11994
rect 21094 11942 21106 11994
rect 21158 11942 23850 11994
rect 23902 11942 23914 11994
rect 23966 11942 23978 11994
rect 24030 11942 24042 11994
rect 24094 11942 24106 11994
rect 24158 11942 24164 11994
rect 1104 11920 24164 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 10597 11883 10655 11889
rect 1627 11852 2774 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 382 11704 388 11756
rect 440 11744 446 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 440 11716 1409 11744
rect 440 11704 446 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 2746 11744 2774 11852
rect 10597 11849 10609 11883
rect 10643 11880 10655 11883
rect 10870 11880 10876 11892
rect 10643 11852 10876 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11204 11852 11529 11880
rect 11204 11840 11210 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11756 11852 11989 11880
rect 11756 11840 11762 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 12529 11883 12587 11889
rect 12529 11880 12541 11883
rect 11977 11843 12035 11849
rect 12084 11852 12541 11880
rect 9214 11812 9220 11824
rect 9140 11784 9220 11812
rect 3234 11744 3240 11756
rect 2746 11716 3240 11744
rect 1397 11707 1455 11713
rect 3234 11704 3240 11716
rect 3292 11744 3298 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 3292 11716 4077 11744
rect 3292 11704 3298 11716
rect 4065 11713 4077 11716
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 4203 11716 4537 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4525 11713 4537 11716
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 5442 11704 5448 11756
rect 5500 11704 5506 11756
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 9140 11753 9168 11784
rect 9214 11772 9220 11784
rect 9272 11812 9278 11824
rect 9582 11812 9588 11824
rect 9272 11784 9588 11812
rect 9272 11772 9278 11784
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 12084 11812 12112 11852
rect 12529 11849 12541 11852
rect 12575 11880 12587 11883
rect 14090 11880 14096 11892
rect 12575 11852 14096 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 16482 11840 16488 11892
rect 16540 11840 16546 11892
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 17678 11880 17684 11892
rect 16991 11852 17684 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18509 11883 18567 11889
rect 18509 11880 18521 11883
rect 18380 11852 18521 11880
rect 18380 11840 18386 11852
rect 18509 11849 18521 11852
rect 18555 11849 18567 11883
rect 18509 11843 18567 11849
rect 19242 11840 19248 11892
rect 19300 11840 19306 11892
rect 20717 11883 20775 11889
rect 20717 11849 20729 11883
rect 20763 11849 20775 11883
rect 20717 11843 20775 11849
rect 13814 11812 13820 11824
rect 10744 11784 12112 11812
rect 12406 11784 13820 11812
rect 10744 11772 10750 11784
rect 9398 11753 9404 11756
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 9392 11744 9404 11753
rect 9359 11716 9404 11744
rect 9125 11707 9183 11713
rect 9392 11707 9404 11716
rect 9398 11704 9404 11707
rect 9456 11704 9462 11756
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10192 11716 10977 11744
rect 10192 11704 10198 11716
rect 10965 11713 10977 11716
rect 11011 11744 11023 11747
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11011 11716 11897 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11885 11713 11897 11716
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 3384 11648 3525 11676
rect 3384 11636 3390 11648
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11676 4399 11679
rect 4890 11676 4896 11688
rect 4387 11648 4896 11676
rect 4387 11645 4399 11648
rect 4341 11639 4399 11645
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5074 11636 5080 11688
rect 5132 11636 5138 11688
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11676 7527 11679
rect 7742 11676 7748 11688
rect 7515 11648 7748 11676
rect 7515 11645 7527 11648
rect 7469 11639 7527 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 8478 11636 8484 11688
rect 8536 11636 8542 11688
rect 11054 11636 11060 11688
rect 11112 11636 11118 11688
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 12161 11679 12219 11685
rect 11204 11648 11560 11676
rect 11204 11636 11210 11648
rect 1670 11568 1676 11620
rect 1728 11608 1734 11620
rect 5261 11611 5319 11617
rect 5261 11608 5273 11611
rect 1728 11580 5273 11608
rect 1728 11568 1734 11580
rect 5261 11577 5273 11580
rect 5307 11577 5319 11611
rect 5261 11571 5319 11577
rect 10505 11611 10563 11617
rect 10505 11577 10517 11611
rect 10551 11608 10563 11611
rect 11422 11608 11428 11620
rect 10551 11580 11428 11608
rect 10551 11577 10563 11580
rect 10505 11571 10563 11577
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 2869 11543 2927 11549
rect 2869 11540 2881 11543
rect 2832 11512 2881 11540
rect 2832 11500 2838 11512
rect 2869 11509 2881 11512
rect 2915 11509 2927 11543
rect 2869 11503 2927 11509
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3697 11543 3755 11549
rect 3697 11540 3709 11543
rect 3476 11512 3709 11540
rect 3476 11500 3482 11512
rect 3697 11509 3709 11512
rect 3743 11509 3755 11543
rect 3697 11503 3755 11509
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 8110 11500 8116 11552
rect 8168 11500 8174 11552
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9398 11540 9404 11552
rect 9079 11512 9404 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 11532 11540 11560 11648
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 12406 11676 12434 11784
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 17402 11821 17408 11824
rect 17396 11812 17408 11821
rect 17363 11784 17408 11812
rect 17396 11775 17408 11784
rect 17402 11772 17408 11775
rect 17460 11772 17466 11824
rect 18690 11772 18696 11824
rect 18748 11812 18754 11824
rect 20732 11812 20760 11843
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21508 11852 21833 11880
rect 21508 11840 21514 11852
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 23474 11812 23480 11824
rect 18748 11784 20760 11812
rect 20916 11784 23480 11812
rect 18748 11772 18754 11784
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 12710 11744 12716 11756
rect 12667 11716 12716 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 12894 11744 12900 11756
rect 12851 11716 12900 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13078 11753 13084 11756
rect 13072 11707 13084 11753
rect 13078 11704 13084 11707
rect 13136 11704 13142 11756
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14240 11716 14657 11744
rect 14240 11704 14246 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14783 11716 15117 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16574 11744 16580 11756
rect 15979 11716 16580 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16761 11747 16819 11753
rect 16761 11713 16773 11747
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 12207 11648 12434 11676
rect 13832 11648 14841 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 13722 11540 13728 11552
rect 11532 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11540 13786 11552
rect 13832 11540 13860 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 14185 11611 14243 11617
rect 14185 11577 14197 11611
rect 14231 11608 14243 11611
rect 15672 11608 15700 11639
rect 15930 11608 15936 11620
rect 14231 11580 15936 11608
rect 14231 11577 14243 11580
rect 14185 11571 14243 11577
rect 15930 11568 15936 11580
rect 15988 11568 15994 11620
rect 16776 11608 16804 11707
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16908 11716 17141 11744
rect 16908 11704 16914 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 18598 11704 18604 11756
rect 18656 11704 18662 11756
rect 20916 11753 20944 11784
rect 23474 11772 23480 11784
rect 23532 11772 23538 11824
rect 20901 11747 20959 11753
rect 20901 11713 20913 11747
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 22327 11716 22753 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22741 11713 22753 11716
rect 22787 11713 22799 11747
rect 22741 11707 22799 11713
rect 23290 11704 23296 11756
rect 23348 11704 23354 11756
rect 23658 11704 23664 11756
rect 23716 11704 23722 11756
rect 21085 11679 21143 11685
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 21174 11676 21180 11688
rect 21131 11648 21180 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 16040 11580 16804 11608
rect 22204 11608 22232 11704
rect 22465 11679 22523 11685
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 22830 11676 22836 11688
rect 22511 11648 22836 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 22830 11636 22836 11648
rect 22888 11636 22894 11688
rect 23477 11611 23535 11617
rect 23477 11608 23489 11611
rect 22204 11580 23489 11608
rect 13780 11512 13860 11540
rect 13780 11500 13786 11512
rect 14274 11500 14280 11552
rect 14332 11500 14338 11552
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 16040 11540 16068 11580
rect 23477 11577 23489 11580
rect 23523 11577 23535 11611
rect 23477 11571 23535 11577
rect 15712 11512 16068 11540
rect 15712 11500 15718 11512
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 21266 11540 21272 11552
rect 16172 11512 21272 11540
rect 16172 11500 16178 11512
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 21634 11500 21640 11552
rect 21692 11500 21698 11552
rect 1104 11450 24012 11472
rect 1104 11398 1350 11450
rect 1402 11398 1414 11450
rect 1466 11398 1478 11450
rect 1530 11398 1542 11450
rect 1594 11398 1606 11450
rect 1658 11398 4350 11450
rect 4402 11398 4414 11450
rect 4466 11398 4478 11450
rect 4530 11398 4542 11450
rect 4594 11398 4606 11450
rect 4658 11398 7350 11450
rect 7402 11398 7414 11450
rect 7466 11398 7478 11450
rect 7530 11398 7542 11450
rect 7594 11398 7606 11450
rect 7658 11398 10350 11450
rect 10402 11398 10414 11450
rect 10466 11398 10478 11450
rect 10530 11398 10542 11450
rect 10594 11398 10606 11450
rect 10658 11398 13350 11450
rect 13402 11398 13414 11450
rect 13466 11398 13478 11450
rect 13530 11398 13542 11450
rect 13594 11398 13606 11450
rect 13658 11398 16350 11450
rect 16402 11398 16414 11450
rect 16466 11398 16478 11450
rect 16530 11398 16542 11450
rect 16594 11398 16606 11450
rect 16658 11398 19350 11450
rect 19402 11398 19414 11450
rect 19466 11398 19478 11450
rect 19530 11398 19542 11450
rect 19594 11398 19606 11450
rect 19658 11398 22350 11450
rect 22402 11398 22414 11450
rect 22466 11398 22478 11450
rect 22530 11398 22542 11450
rect 22594 11398 22606 11450
rect 22658 11398 24012 11450
rect 1104 11376 24012 11398
rect 8110 11336 8116 11348
rect 2056 11308 8116 11336
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 2056 11141 2084 11308
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 8720 11308 9965 11336
rect 8720 11296 8726 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 9953 11299 10011 11305
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11112 11308 11805 11336
rect 11112 11296 11118 11308
rect 11793 11305 11805 11308
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13078 11336 13084 11348
rect 13035 11308 13084 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13722 11336 13728 11348
rect 13403 11308 13728 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 13872 11308 14197 11336
rect 13872 11296 13878 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14185 11299 14243 11305
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 16114 11336 16120 11348
rect 15335 11308 16120 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11336 17279 11339
rect 17494 11336 17500 11348
rect 17267 11308 17500 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18690 11336 18696 11348
rect 17604 11308 18696 11336
rect 2409 11271 2467 11277
rect 2409 11237 2421 11271
rect 2455 11237 2467 11271
rect 2409 11231 2467 11237
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2424 11132 2452 11231
rect 3602 11228 3608 11280
rect 3660 11228 3666 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 13004 11240 13645 11268
rect 13004 11212 13032 11240
rect 13633 11237 13645 11240
rect 13679 11268 13691 11271
rect 15470 11268 15476 11280
rect 13679 11240 15476 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3510 11200 3516 11212
rect 3099 11172 3516 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 3510 11160 3516 11172
rect 3568 11200 3574 11212
rect 3694 11200 3700 11212
rect 3568 11172 3700 11200
rect 3568 11160 3574 11172
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10686 11200 10692 11212
rect 10643 11172 10692 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11422 11160 11428 11212
rect 11480 11160 11486 11212
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 12526 11200 12532 11212
rect 12483 11172 12532 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12986 11160 12992 11212
rect 13044 11160 13050 11212
rect 14274 11200 14280 11212
rect 13188 11172 14280 11200
rect 2363 11104 2452 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 3786 11092 3792 11144
rect 3844 11141 3850 11144
rect 3844 11132 3854 11141
rect 3844 11104 3889 11132
rect 3844 11095 3854 11104
rect 3844 11092 3850 11095
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5408 11104 5457 11132
rect 5408 11092 5414 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 6963 11104 8493 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 8481 11101 8493 11104
rect 8527 11132 8539 11135
rect 8527 11104 9628 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9600 11076 9628 11104
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 13188 11141 13216 11172
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 10192 11104 10333 11132
rect 10192 11092 10198 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 15120 11141 15148 11240
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 16577 11271 16635 11277
rect 16577 11237 16589 11271
rect 16623 11268 16635 11271
rect 17310 11268 17316 11280
rect 16623 11240 17316 11268
rect 16623 11237 16635 11240
rect 16577 11231 16635 11237
rect 17310 11228 17316 11240
rect 17368 11228 17374 11280
rect 17604 11141 17632 11308
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 21818 11336 21824 11348
rect 21131 11308 21824 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 21818 11296 21824 11308
rect 21876 11336 21882 11348
rect 21876 11308 23428 11336
rect 21876 11296 21882 11308
rect 20714 11228 20720 11280
rect 20772 11268 20778 11280
rect 21177 11271 21235 11277
rect 21177 11268 21189 11271
rect 20772 11240 21189 11268
rect 20772 11228 20778 11240
rect 21177 11237 21189 11240
rect 21223 11237 21235 11271
rect 21177 11231 21235 11237
rect 21450 11228 21456 11280
rect 21508 11268 21514 11280
rect 22005 11271 22063 11277
rect 22005 11268 22017 11271
rect 21508 11240 22017 11268
rect 21508 11228 21514 11240
rect 22005 11237 22017 11240
rect 22051 11237 22063 11271
rect 22005 11231 22063 11237
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13320 11104 13461 11132
rect 13320 11092 13326 11104
rect 13449 11101 13461 11104
rect 13495 11132 13507 11135
rect 15105 11135 15163 11141
rect 13495 11104 14780 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 3234 11064 3240 11076
rect 2915 11036 3240 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 4034 11067 4092 11073
rect 4034 11064 4046 11067
rect 3660 11036 4046 11064
rect 3660 11024 3666 11036
rect 4034 11033 4046 11036
rect 4080 11033 4092 11067
rect 4034 11027 4092 11033
rect 5712 11067 5770 11073
rect 5712 11033 5724 11067
rect 5758 11064 5770 11067
rect 6454 11064 6460 11076
rect 5758 11036 6460 11064
rect 5758 11033 5770 11036
rect 5712 11027 5770 11033
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7162 11067 7220 11073
rect 7162 11064 7174 11067
rect 7064 11036 7174 11064
rect 7064 11024 7070 11036
rect 7162 11033 7174 11036
rect 7208 11033 7220 11067
rect 7162 11027 7220 11033
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 8938 11064 8944 11076
rect 8260 11036 8944 11064
rect 8260 11024 8266 11036
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 9677 11067 9735 11073
rect 9677 11064 9689 11067
rect 9640 11036 9689 11064
rect 9640 11024 9646 11036
rect 9677 11033 9689 11036
rect 9723 11033 9735 11067
rect 9677 11027 9735 11033
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11064 10471 11067
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 10459 11036 10793 11064
rect 10459 11033 10471 11036
rect 10413 11027 10471 11033
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 10781 11027 10839 11033
rect 13817 11067 13875 11073
rect 13817 11033 13829 11067
rect 13863 11064 13875 11067
rect 13998 11064 14004 11076
rect 13863 11036 14004 11064
rect 13863 11033 13875 11036
rect 13817 11027 13875 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14274 11024 14280 11076
rect 14332 11024 14338 11076
rect 14752 11064 14780 11104
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11101 17647 11135
rect 17880 11132 17908 11163
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18693 11203 18751 11209
rect 18693 11200 18705 11203
rect 18380 11172 18705 11200
rect 18380 11160 18386 11172
rect 18693 11169 18705 11172
rect 18739 11169 18751 11203
rect 18693 11163 18751 11169
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 23400 11209 23428 11308
rect 21729 11203 21787 11209
rect 21729 11200 21741 11203
rect 21324 11172 21741 11200
rect 21324 11160 21330 11172
rect 21729 11169 21741 11172
rect 21775 11169 21787 11203
rect 22557 11203 22615 11209
rect 22557 11200 22569 11203
rect 21729 11163 21787 11169
rect 21836 11172 22569 11200
rect 19705 11135 19763 11141
rect 17880 11104 18368 11132
rect 17589 11095 17647 11101
rect 15654 11064 15660 11076
rect 14752 11036 15660 11064
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 16390 11024 16396 11076
rect 16448 11024 16454 11076
rect 17681 11067 17739 11073
rect 17681 11033 17693 11067
rect 17727 11064 17739 11067
rect 18141 11067 18199 11073
rect 18141 11064 18153 11067
rect 17727 11036 18153 11064
rect 17727 11033 17739 11036
rect 17681 11027 17739 11033
rect 18141 11033 18153 11036
rect 18187 11033 18199 11067
rect 18340 11064 18368 11104
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 19794 11132 19800 11144
rect 19751 11104 19800 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 20438 11132 20444 11144
rect 19904 11104 20444 11132
rect 19904 11064 19932 11104
rect 20438 11092 20444 11104
rect 20496 11132 20502 11144
rect 21836 11132 21864 11172
rect 22557 11169 22569 11172
rect 22603 11169 22615 11203
rect 22557 11163 22615 11169
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11169 23443 11203
rect 23385 11163 23443 11169
rect 20496 11104 21864 11132
rect 20496 11092 20502 11104
rect 22002 11092 22008 11144
rect 22060 11132 22066 11144
rect 22373 11135 22431 11141
rect 22373 11132 22385 11135
rect 22060 11104 22385 11132
rect 22060 11092 22066 11104
rect 22373 11101 22385 11104
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 18340 11036 19932 11064
rect 19972 11067 20030 11073
rect 18141 11027 18199 11033
rect 19972 11033 19984 11067
rect 20018 11064 20030 11067
rect 20070 11064 20076 11076
rect 20018 11036 20076 11064
rect 20018 11033 20030 11036
rect 19972 11027 20030 11033
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 21545 11067 21603 11073
rect 21545 11033 21557 11067
rect 21591 11064 21603 11067
rect 22833 11067 22891 11073
rect 22833 11064 22845 11067
rect 21591 11036 21864 11064
rect 21591 11033 21603 11036
rect 21545 11027 21603 11033
rect 1486 10956 1492 11008
rect 1544 10956 1550 11008
rect 1854 10956 1860 11008
rect 1912 10956 1918 11008
rect 2130 10956 2136 11008
rect 2188 10956 2194 11008
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 4246 10996 4252 11008
rect 3384 10968 4252 10996
rect 3384 10956 3390 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5169 10999 5227 11005
rect 5169 10996 5181 10999
rect 5132 10968 5181 10996
rect 5132 10956 5138 10968
rect 5169 10965 5181 10968
rect 5215 10965 5227 10999
rect 5169 10959 5227 10965
rect 6825 10999 6883 11005
rect 6825 10965 6837 10999
rect 6871 10996 6883 10999
rect 7742 10996 7748 11008
rect 6871 10968 7748 10996
rect 6871 10965 6883 10968
rect 6825 10959 6883 10965
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 8478 10996 8484 11008
rect 8343 10968 8484 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 21266 10956 21272 11008
rect 21324 10996 21330 11008
rect 21637 10999 21695 11005
rect 21637 10996 21649 10999
rect 21324 10968 21649 10996
rect 21324 10956 21330 10968
rect 21637 10965 21649 10968
rect 21683 10965 21695 10999
rect 21836 10996 21864 11036
rect 22204 11036 22845 11064
rect 22204 10996 22232 11036
rect 22833 11033 22845 11036
rect 22879 11033 22891 11067
rect 22833 11027 22891 11033
rect 21836 10968 22232 10996
rect 22465 10999 22523 11005
rect 21637 10959 21695 10965
rect 22465 10965 22477 10999
rect 22511 10996 22523 10999
rect 23014 10996 23020 11008
rect 22511 10968 23020 10996
rect 22511 10965 22523 10968
rect 22465 10959 22523 10965
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 1104 10906 24164 10928
rect 1104 10854 2850 10906
rect 2902 10854 2914 10906
rect 2966 10854 2978 10906
rect 3030 10854 3042 10906
rect 3094 10854 3106 10906
rect 3158 10854 5850 10906
rect 5902 10854 5914 10906
rect 5966 10854 5978 10906
rect 6030 10854 6042 10906
rect 6094 10854 6106 10906
rect 6158 10854 8850 10906
rect 8902 10854 8914 10906
rect 8966 10854 8978 10906
rect 9030 10854 9042 10906
rect 9094 10854 9106 10906
rect 9158 10854 11850 10906
rect 11902 10854 11914 10906
rect 11966 10854 11978 10906
rect 12030 10854 12042 10906
rect 12094 10854 12106 10906
rect 12158 10854 14850 10906
rect 14902 10854 14914 10906
rect 14966 10854 14978 10906
rect 15030 10854 15042 10906
rect 15094 10854 15106 10906
rect 15158 10854 17850 10906
rect 17902 10854 17914 10906
rect 17966 10854 17978 10906
rect 18030 10854 18042 10906
rect 18094 10854 18106 10906
rect 18158 10854 20850 10906
rect 20902 10854 20914 10906
rect 20966 10854 20978 10906
rect 21030 10854 21042 10906
rect 21094 10854 21106 10906
rect 21158 10854 23850 10906
rect 23902 10854 23914 10906
rect 23966 10854 23978 10906
rect 24030 10854 24042 10906
rect 24094 10854 24106 10906
rect 24158 10854 24164 10906
rect 1104 10832 24164 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3326 10792 3332 10804
rect 2915 10764 3332 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 5074 10792 5080 10804
rect 3528 10764 5080 10792
rect 1756 10727 1814 10733
rect 1756 10693 1768 10727
rect 1802 10724 1814 10727
rect 2130 10724 2136 10736
rect 1802 10696 2136 10724
rect 1802 10693 1814 10696
rect 1756 10687 1814 10693
rect 2130 10684 2136 10696
rect 2188 10684 2194 10736
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3418 10656 3424 10668
rect 3099 10628 3424 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 3528 10656 3556 10764
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5442 10792 5448 10804
rect 5215 10764 5448 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6917 10795 6975 10801
rect 6917 10761 6929 10795
rect 6963 10792 6975 10795
rect 7006 10792 7012 10804
rect 6963 10764 7012 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 7116 10764 8953 10792
rect 6178 10684 6184 10736
rect 6236 10684 6242 10736
rect 3528 10628 3648 10656
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10557 1547 10591
rect 1489 10551 1547 10557
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 1504 10452 1532 10551
rect 3344 10520 3372 10551
rect 3510 10548 3516 10600
rect 3568 10548 3574 10600
rect 3620 10520 3648 10628
rect 4246 10616 4252 10668
rect 4304 10616 4310 10668
rect 6362 10616 6368 10668
rect 6420 10616 6426 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7116 10656 7144 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 9398 10752 9404 10804
rect 9456 10752 9462 10804
rect 20809 10795 20867 10801
rect 20809 10761 20821 10795
rect 20855 10792 20867 10795
rect 21174 10792 21180 10804
rect 20855 10764 21180 10792
rect 20855 10761 20867 10764
rect 20809 10755 20867 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 21361 10795 21419 10801
rect 21361 10761 21373 10795
rect 21407 10792 21419 10795
rect 21634 10792 21640 10804
rect 21407 10764 21640 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 22097 10795 22155 10801
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 23382 10792 23388 10804
rect 22143 10764 23388 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12805 10727 12863 10733
rect 12805 10724 12817 10727
rect 12032 10696 12817 10724
rect 12032 10684 12038 10696
rect 12805 10693 12817 10696
rect 12851 10724 12863 10727
rect 16117 10727 16175 10733
rect 16117 10724 16129 10727
rect 12851 10696 16129 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 16117 10693 16129 10696
rect 16163 10724 16175 10727
rect 16390 10724 16396 10736
rect 16163 10696 16396 10724
rect 16163 10693 16175 10696
rect 16117 10687 16175 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 21266 10684 21272 10736
rect 21324 10724 21330 10736
rect 22002 10724 22008 10736
rect 21324 10696 22008 10724
rect 21324 10684 21330 10696
rect 22002 10684 22008 10696
rect 22060 10684 22066 10736
rect 6779 10628 7144 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7650 10616 7656 10668
rect 7708 10616 7714 10668
rect 7742 10616 7748 10668
rect 7800 10665 7806 10668
rect 7800 10659 7849 10665
rect 7800 10625 7803 10659
rect 7837 10625 7849 10659
rect 7800 10619 7849 10625
rect 7800 10616 7806 10619
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 8849 10659 8907 10665
rect 8849 10656 8861 10659
rect 8536 10628 8861 10656
rect 8536 10616 8542 10628
rect 8849 10625 8861 10628
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 11238 10656 11244 10668
rect 9999 10628 11244 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 11238 10616 11244 10628
rect 11296 10656 11302 10668
rect 11296 10628 12434 10656
rect 11296 10616 11302 10628
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 4366 10591 4424 10597
rect 4366 10588 4378 10591
rect 3936 10560 4378 10588
rect 3936 10548 3942 10560
rect 4366 10557 4378 10560
rect 4412 10557 4424 10591
rect 4366 10551 4424 10557
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4706 10588 4712 10600
rect 4571 10560 4712 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4706 10548 4712 10560
rect 4764 10588 4770 10600
rect 4890 10588 4896 10600
rect 4764 10560 4896 10588
rect 4764 10548 4770 10560
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 5626 10548 5632 10600
rect 5684 10588 5690 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 5684 10560 7941 10588
rect 5684 10548 5690 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 8570 10588 8576 10600
rect 8251 10560 8576 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 8754 10588 8760 10600
rect 8711 10560 8760 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9456 10560 9505 10588
rect 9456 10548 9462 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 3344 10492 3648 10520
rect 3973 10523 4031 10529
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4062 10520 4068 10532
rect 4019 10492 4068 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 4908 10520 4936 10548
rect 7190 10520 7196 10532
rect 4908 10492 7196 10520
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 12406 10520 12434 10628
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 19702 10665 19708 10668
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14148 10628 14841 10656
rect 14148 10616 14154 10628
rect 14829 10625 14841 10628
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 19696 10619 19708 10665
rect 19702 10616 19708 10619
rect 19760 10616 19766 10668
rect 21910 10616 21916 10668
rect 21968 10616 21974 10668
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22445 10659 22503 10665
rect 22445 10656 22457 10659
rect 22152 10628 22457 10656
rect 22152 10616 22158 10628
rect 22445 10625 22457 10628
rect 22491 10625 22503 10659
rect 22445 10619 22503 10625
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 15068 10560 15117 10588
rect 15068 10548 15074 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16669 10591 16727 10597
rect 16669 10588 16681 10591
rect 15896 10560 16681 10588
rect 15896 10548 15902 10560
rect 16669 10557 16681 10560
rect 16715 10557 16727 10591
rect 16669 10551 16727 10557
rect 19429 10591 19487 10597
rect 19429 10557 19441 10591
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10588 21603 10591
rect 21726 10588 21732 10600
rect 21591 10560 21732 10588
rect 21591 10557 21603 10560
rect 21545 10551 21603 10557
rect 12618 10520 12624 10532
rect 12406 10492 12624 10520
rect 12618 10480 12624 10492
rect 12676 10520 12682 10532
rect 12986 10520 12992 10532
rect 12676 10492 12992 10520
rect 12676 10480 12682 10492
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 1854 10452 1860 10464
rect 1504 10424 1860 10452
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 4890 10452 4896 10464
rect 3283 10424 4896 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6730 10452 6736 10464
rect 6595 10424 6736 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 8294 10452 8300 10464
rect 7055 10424 8300 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 8720 10424 9873 10452
rect 8720 10412 8726 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14516 10424 15025 10452
rect 14516 10412 14522 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 15746 10412 15752 10464
rect 15804 10412 15810 10464
rect 16025 10455 16083 10461
rect 16025 10421 16037 10455
rect 16071 10452 16083 10455
rect 16206 10452 16212 10464
rect 16071 10424 16212 10452
rect 16071 10421 16083 10424
rect 16025 10415 16083 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 17310 10412 17316 10464
rect 17368 10412 17374 10464
rect 19444 10452 19472 10551
rect 21726 10548 21732 10560
rect 21784 10548 21790 10600
rect 22189 10591 22247 10597
rect 22189 10557 22201 10591
rect 22235 10557 22247 10591
rect 22189 10551 22247 10557
rect 22204 10520 22232 10551
rect 20364 10492 22232 10520
rect 19794 10452 19800 10464
rect 19444 10424 19800 10452
rect 19794 10412 19800 10424
rect 19852 10452 19858 10464
rect 20364 10452 20392 10492
rect 19852 10424 20392 10452
rect 19852 10412 19858 10424
rect 20898 10412 20904 10464
rect 20956 10412 20962 10464
rect 23566 10412 23572 10464
rect 23624 10412 23630 10464
rect 1104 10362 24012 10384
rect 1104 10310 1350 10362
rect 1402 10310 1414 10362
rect 1466 10310 1478 10362
rect 1530 10310 1542 10362
rect 1594 10310 1606 10362
rect 1658 10310 4350 10362
rect 4402 10310 4414 10362
rect 4466 10310 4478 10362
rect 4530 10310 4542 10362
rect 4594 10310 4606 10362
rect 4658 10310 7350 10362
rect 7402 10310 7414 10362
rect 7466 10310 7478 10362
rect 7530 10310 7542 10362
rect 7594 10310 7606 10362
rect 7658 10310 10350 10362
rect 10402 10310 10414 10362
rect 10466 10310 10478 10362
rect 10530 10310 10542 10362
rect 10594 10310 10606 10362
rect 10658 10310 13350 10362
rect 13402 10310 13414 10362
rect 13466 10310 13478 10362
rect 13530 10310 13542 10362
rect 13594 10310 13606 10362
rect 13658 10310 16350 10362
rect 16402 10310 16414 10362
rect 16466 10310 16478 10362
rect 16530 10310 16542 10362
rect 16594 10310 16606 10362
rect 16658 10310 19350 10362
rect 19402 10310 19414 10362
rect 19466 10310 19478 10362
rect 19530 10310 19542 10362
rect 19594 10310 19606 10362
rect 19658 10310 22350 10362
rect 22402 10310 22414 10362
rect 22466 10310 22478 10362
rect 22530 10310 22542 10362
rect 22594 10310 22606 10362
rect 22658 10310 24012 10362
rect 1104 10288 24012 10310
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4798 10248 4804 10260
rect 4212 10220 4804 10248
rect 4212 10208 4218 10220
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5626 10208 5632 10260
rect 5684 10208 5690 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8662 10248 8668 10260
rect 7800 10220 8668 10248
rect 7800 10208 7806 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 8754 10208 8760 10260
rect 8812 10208 8818 10260
rect 11974 10208 11980 10260
rect 12032 10208 12038 10260
rect 14090 10208 14096 10260
rect 14148 10208 14154 10260
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19760 10220 19809 10248
rect 19760 10208 19766 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 19797 10211 19855 10217
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 21324 10220 21956 10248
rect 21324 10208 21330 10220
rect 3510 10180 3516 10192
rect 3068 10152 3516 10180
rect 3068 10121 3096 10152
rect 3510 10140 3516 10152
rect 3568 10180 3574 10192
rect 3789 10183 3847 10189
rect 3789 10180 3801 10183
rect 3568 10152 3801 10180
rect 3568 10140 3574 10152
rect 3789 10149 3801 10152
rect 3835 10149 3847 10183
rect 3789 10143 3847 10149
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10081 3111 10115
rect 3053 10075 3111 10081
rect 3605 10115 3663 10121
rect 3605 10081 3617 10115
rect 3651 10112 3663 10115
rect 4154 10112 4160 10124
rect 3651 10084 4160 10112
rect 3651 10081 3663 10084
rect 3605 10075 3663 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 8772 10112 8800 10208
rect 12986 10140 12992 10192
rect 13044 10180 13050 10192
rect 13044 10152 13860 10180
rect 13044 10140 13050 10152
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 7055 10084 7420 10112
rect 8772 10084 9505 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 3786 10044 3792 10056
rect 1535 10016 1900 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 1872 9988 1900 10016
rect 2746 10016 3792 10044
rect 1762 9985 1768 9988
rect 1756 9939 1768 9985
rect 1762 9936 1768 9939
rect 1820 9936 1826 9988
rect 1854 9936 1860 9988
rect 1912 9976 1918 9988
rect 2746 9976 2774 10016
rect 3786 10004 3792 10016
rect 3844 10044 3850 10056
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 3844 10016 5181 10044
rect 3844 10004 3850 10016
rect 5169 10013 5181 10016
rect 5215 10044 5227 10047
rect 5350 10044 5356 10056
rect 5215 10016 5356 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 6730 10004 6736 10056
rect 6788 10053 6794 10056
rect 6788 10044 6800 10053
rect 6788 10016 6833 10044
rect 6788 10007 6800 10016
rect 6788 10004 6794 10007
rect 7098 10004 7104 10056
rect 7156 10004 7162 10056
rect 7392 10053 7420 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 9640 10084 10241 10112
rect 9640 10072 9646 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 13722 10072 13728 10124
rect 13780 10072 13786 10124
rect 13832 10112 13860 10152
rect 15286 10140 15292 10192
rect 15344 10140 15350 10192
rect 17773 10183 17831 10189
rect 17773 10149 17785 10183
rect 17819 10180 17831 10183
rect 17819 10152 18460 10180
rect 17819 10149 17831 10152
rect 17773 10143 17831 10149
rect 13832 10084 14780 10112
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7423 10016 8340 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 8312 9988 8340 10016
rect 13170 10004 13176 10056
rect 13228 10004 13234 10056
rect 14752 10053 14780 10084
rect 15010 10072 15016 10124
rect 15068 10072 15074 10124
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10112 15807 10115
rect 15838 10112 15844 10124
rect 15795 10084 15844 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 15930 10072 15936 10124
rect 15988 10072 15994 10124
rect 18432 10121 18460 10152
rect 20898 10140 20904 10192
rect 20956 10140 20962 10192
rect 21928 10189 21956 10220
rect 23014 10208 23020 10260
rect 23072 10208 23078 10260
rect 21913 10183 21971 10189
rect 21913 10149 21925 10183
rect 21959 10149 21971 10183
rect 21913 10143 21971 10149
rect 18417 10115 18475 10121
rect 18417 10081 18429 10115
rect 18463 10112 18475 10115
rect 18506 10112 18512 10124
rect 18463 10084 18512 10112
rect 18463 10081 18475 10084
rect 18417 10075 18475 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 20916 10112 20944 10140
rect 19996 10084 20944 10112
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 14737 10047 14795 10053
rect 13587 10016 14228 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 1912 9948 2774 9976
rect 1912 9936 1918 9948
rect 4890 9936 4896 9988
rect 4948 9985 4954 9988
rect 4948 9976 4960 9985
rect 7622 9979 7680 9985
rect 7622 9976 7634 9979
rect 4948 9948 4993 9976
rect 7300 9948 7634 9976
rect 4948 9939 4960 9948
rect 4948 9936 4954 9939
rect 2869 9911 2927 9917
rect 2869 9877 2881 9911
rect 2915 9908 2927 9911
rect 3878 9908 3884 9920
rect 2915 9880 3884 9908
rect 2915 9877 2927 9880
rect 2869 9871 2927 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 7300 9917 7328 9948
rect 7622 9945 7634 9948
rect 7668 9945 7680 9979
rect 7622 9939 7680 9945
rect 8294 9936 8300 9988
rect 8352 9936 8358 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8444 9948 8953 9976
rect 8444 9936 8450 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 10502 9936 10508 9988
rect 10560 9936 10566 9988
rect 11054 9936 11060 9988
rect 11112 9936 11118 9988
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 13188 9976 13216 10004
rect 14200 9988 14228 10016
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 14826 10004 14832 10056
rect 14884 10053 14890 10056
rect 14884 10047 14933 10053
rect 14884 10013 14887 10047
rect 14921 10013 14933 10047
rect 14884 10007 14933 10013
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 14884 10004 14890 10007
rect 12492 9948 13952 9976
rect 12492 9936 12498 9948
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 12584 9880 13185 9908
rect 12584 9868 12590 9880
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 13173 9871 13231 9877
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 13814 9908 13820 9920
rect 13679 9880 13820 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 13924 9908 13952 9948
rect 14182 9936 14188 9988
rect 14240 9936 14246 9988
rect 16040 9908 16068 10007
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 19996 10053 20024 10084
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 21499 10115 21557 10121
rect 21499 10112 21511 10115
rect 21232 10084 21511 10112
rect 21232 10072 21238 10084
rect 21499 10081 21511 10084
rect 21545 10081 21557 10115
rect 21499 10075 21557 10081
rect 21637 10115 21695 10121
rect 21637 10081 21649 10115
rect 21683 10112 21695 10115
rect 21818 10112 21824 10124
rect 21683 10084 21824 10112
rect 21683 10081 21695 10084
rect 21637 10075 21695 10081
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 22373 10115 22431 10121
rect 22373 10081 22385 10115
rect 22419 10112 22431 10115
rect 23566 10112 23572 10124
rect 22419 10084 23572 10112
rect 22419 10081 22431 10084
rect 22373 10075 22431 10081
rect 23566 10072 23572 10084
rect 23624 10072 23630 10124
rect 16393 10047 16451 10053
rect 16393 10044 16405 10047
rect 16172 10016 16405 10044
rect 16172 10004 16178 10016
rect 16393 10013 16405 10016
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10044 20315 10047
rect 20714 10044 20720 10056
rect 20303 10016 20720 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 21358 10004 21364 10056
rect 21416 10004 21422 10056
rect 22186 10004 22192 10056
rect 22244 10044 22250 10056
rect 22557 10047 22615 10053
rect 22557 10044 22569 10047
rect 22244 10016 22569 10044
rect 22244 10004 22250 10016
rect 22557 10013 22569 10016
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 16666 9985 16672 9988
rect 16660 9939 16672 9985
rect 16666 9936 16672 9939
rect 16724 9936 16730 9988
rect 13924 9880 16068 9908
rect 16206 9868 16212 9920
rect 16264 9868 16270 9920
rect 17126 9868 17132 9920
rect 17184 9908 17190 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17184 9880 17877 9908
rect 17184 9868 17190 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 20717 9911 20775 9917
rect 20717 9877 20729 9911
rect 20763 9908 20775 9911
rect 22738 9908 22744 9920
rect 20763 9880 22744 9908
rect 20763 9877 20775 9880
rect 20717 9871 20775 9877
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 22830 9868 22836 9920
rect 22888 9868 22894 9920
rect 1104 9818 24164 9840
rect 1104 9766 2850 9818
rect 2902 9766 2914 9818
rect 2966 9766 2978 9818
rect 3030 9766 3042 9818
rect 3094 9766 3106 9818
rect 3158 9766 5850 9818
rect 5902 9766 5914 9818
rect 5966 9766 5978 9818
rect 6030 9766 6042 9818
rect 6094 9766 6106 9818
rect 6158 9766 8850 9818
rect 8902 9766 8914 9818
rect 8966 9766 8978 9818
rect 9030 9766 9042 9818
rect 9094 9766 9106 9818
rect 9158 9766 11850 9818
rect 11902 9766 11914 9818
rect 11966 9766 11978 9818
rect 12030 9766 12042 9818
rect 12094 9766 12106 9818
rect 12158 9766 14850 9818
rect 14902 9766 14914 9818
rect 14966 9766 14978 9818
rect 15030 9766 15042 9818
rect 15094 9766 15106 9818
rect 15158 9766 17850 9818
rect 17902 9766 17914 9818
rect 17966 9766 17978 9818
rect 18030 9766 18042 9818
rect 18094 9766 18106 9818
rect 18158 9766 20850 9818
rect 20902 9766 20914 9818
rect 20966 9766 20978 9818
rect 21030 9766 21042 9818
rect 21094 9766 21106 9818
rect 21158 9766 23850 9818
rect 23902 9766 23914 9818
rect 23966 9766 23978 9818
rect 24030 9766 24042 9818
rect 24094 9766 24106 9818
rect 24158 9766 24164 9818
rect 1104 9744 24164 9766
rect 1762 9664 1768 9716
rect 1820 9704 1826 9716
rect 1949 9707 2007 9713
rect 1949 9704 1961 9707
rect 1820 9676 1961 9704
rect 1820 9664 1826 9676
rect 1949 9673 1961 9676
rect 1995 9673 2007 9707
rect 1949 9667 2007 9673
rect 3234 9664 3240 9716
rect 3292 9664 3298 9716
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 4065 9707 4123 9713
rect 4065 9704 4077 9707
rect 3476 9676 4077 9704
rect 3476 9664 3482 9676
rect 4065 9673 4077 9676
rect 4111 9673 4123 9707
rect 4065 9667 4123 9673
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6362 9704 6368 9716
rect 6227 9676 6368 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7377 9707 7435 9713
rect 7377 9704 7389 9707
rect 7156 9676 7389 9704
rect 7156 9664 7162 9676
rect 7377 9673 7389 9676
rect 7423 9673 7435 9707
rect 9306 9704 9312 9716
rect 7377 9667 7435 9673
rect 8128 9676 9312 9704
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 3252 9636 3280 9664
rect 2823 9608 4016 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 382 9528 388 9580
rect 440 9568 446 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 440 9540 1409 9568
rect 440 9528 446 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 2869 9571 2927 9577
rect 2179 9540 2452 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 2424 9441 2452 9540
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 2915 9540 3249 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3878 9528 3884 9580
rect 3936 9528 3942 9580
rect 3988 9568 4016 9608
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 4212 9608 4537 9636
rect 4212 9596 4218 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 6638 9636 6644 9648
rect 4525 9599 4583 9605
rect 4632 9608 6644 9636
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 3988 9540 4445 9568
rect 4433 9537 4445 9540
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9401 2467 9435
rect 2409 9395 2467 9401
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 3068 9432 3096 9463
rect 4632 9432 4660 9608
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 6822 9596 6828 9648
rect 6880 9596 6886 9648
rect 8128 9636 8156 9676
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10502 9664 10508 9716
rect 10560 9664 10566 9716
rect 14277 9707 14335 9713
rect 14277 9673 14289 9707
rect 14323 9704 14335 9707
rect 14550 9704 14556 9716
rect 14323 9676 14556 9704
rect 14323 9673 14335 9676
rect 14277 9667 14335 9673
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9673 15439 9707
rect 15381 9667 15439 9673
rect 7760 9608 8156 9636
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 7760 9577 7788 9608
rect 8202 9596 8208 9648
rect 8260 9596 8266 9648
rect 9214 9596 9220 9648
rect 9272 9636 9278 9648
rect 15396 9636 15424 9667
rect 15746 9664 15752 9716
rect 15804 9664 15810 9716
rect 16485 9707 16543 9713
rect 16485 9673 16497 9707
rect 16531 9704 16543 9707
rect 16666 9704 16672 9716
rect 16531 9676 16672 9704
rect 16531 9673 16543 9676
rect 16485 9667 16543 9673
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 17129 9707 17187 9713
rect 17129 9673 17141 9707
rect 17175 9704 17187 9707
rect 17310 9704 17316 9716
rect 17175 9676 17316 9704
rect 17175 9673 17187 9676
rect 17129 9667 17187 9673
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 20809 9707 20867 9713
rect 20809 9673 20821 9707
rect 20855 9673 20867 9707
rect 20809 9667 20867 9673
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 9272 9608 10640 9636
rect 9272 9596 9278 9608
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 6779 9540 7757 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8386 9568 8392 9580
rect 7883 9540 8392 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 5258 9500 5264 9512
rect 4755 9472 5264 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5534 9460 5540 9512
rect 5592 9460 5598 9512
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 5644 9472 5733 9500
rect 2832 9404 4660 9432
rect 2832 9392 2838 9404
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 5644 9364 5672 9472
rect 5721 9469 5733 9472
rect 5767 9500 5779 9503
rect 6748 9500 6776 9531
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10612 9577 10640 9608
rect 12636 9608 15424 9636
rect 15856 9608 17049 9636
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9537 10655 9571
rect 10597 9531 10655 9537
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 12526 9568 12532 9580
rect 12391 9540 12532 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 5767 9472 6776 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6880 9472 6929 9500
rect 6880 9460 6886 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7926 9460 7932 9512
rect 7984 9460 7990 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9490 9500 9496 9512
rect 9079 9472 9496 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10428 9500 10456 9531
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12636 9577 12664 9608
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 13153 9571 13211 9577
rect 13153 9568 13165 9571
rect 13004 9540 13165 9568
rect 13004 9500 13032 9540
rect 13153 9537 13165 9540
rect 13199 9537 13211 9571
rect 13153 9531 13211 9537
rect 14366 9528 14372 9580
rect 14424 9528 14430 9580
rect 15856 9577 15884 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 20824 9636 20852 9667
rect 22646 9664 22652 9716
rect 22704 9664 22710 9716
rect 22664 9636 22692 9664
rect 17037 9599 17095 9605
rect 19720 9608 20668 9636
rect 20824 9608 22692 9636
rect 15841 9571 15899 9577
rect 15841 9568 15853 9571
rect 15120 9540 15853 9568
rect 9732 9472 10456 9500
rect 12820 9472 13032 9500
rect 9732 9460 9738 9472
rect 12820 9441 12848 9472
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 15120 9500 15148 9540
rect 15841 9537 15853 9540
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16758 9568 16764 9580
rect 16347 9540 16764 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 18506 9528 18512 9580
rect 18564 9528 18570 9580
rect 19720 9568 19748 9608
rect 19168 9540 19748 9568
rect 14240 9472 15148 9500
rect 14240 9460 14246 9472
rect 15194 9460 15200 9512
rect 15252 9460 15258 9512
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 15948 9432 15976 9463
rect 17218 9460 17224 9512
rect 17276 9460 17282 9512
rect 18230 9500 18236 9512
rect 17880 9472 18236 9500
rect 14608 9404 15976 9432
rect 14608 9392 14614 9404
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 17880 9432 17908 9472
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18414 9509 18420 9512
rect 18392 9503 18420 9509
rect 18392 9469 18404 9503
rect 18392 9463 18420 9469
rect 18414 9460 18420 9463
rect 18472 9460 18478 9512
rect 19168 9500 19196 9540
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 20640 9577 20668 9608
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19852 9540 20269 9568
rect 19852 9528 19858 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 21315 9540 21404 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 18708 9472 19196 9500
rect 16356 9404 17908 9432
rect 16356 9392 16362 9404
rect 1627 9336 5672 9364
rect 6365 9367 6423 9373
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6638 9364 6644 9376
rect 6411 9336 6644 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 10778 9364 10784 9376
rect 10367 9336 10784 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12529 9367 12587 9373
rect 12529 9333 12541 9367
rect 12575 9364 12587 9367
rect 12618 9364 12624 9376
rect 12575 9336 12624 9364
rect 12575 9333 12587 9336
rect 12529 9327 12587 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 15344 9336 16681 9364
rect 15344 9324 15350 9336
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 16669 9327 16727 9333
rect 17589 9367 17647 9373
rect 17589 9333 17601 9367
rect 17635 9364 17647 9367
rect 18708 9364 18736 9472
rect 19242 9460 19248 9512
rect 19300 9460 19306 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19475 9472 20085 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 18785 9435 18843 9441
rect 18785 9401 18797 9435
rect 18831 9432 18843 9435
rect 19058 9432 19064 9444
rect 18831 9404 19064 9432
rect 18831 9401 18843 9404
rect 18785 9395 18843 9401
rect 19058 9392 19064 9404
rect 19116 9392 19122 9444
rect 19150 9392 19156 9444
rect 19208 9432 19214 9444
rect 19444 9432 19472 9463
rect 19208 9404 19472 9432
rect 19208 9392 19214 9404
rect 19610 9392 19616 9444
rect 19668 9432 19674 9444
rect 20438 9432 20444 9444
rect 19668 9404 20444 9432
rect 19668 9392 19674 9404
rect 20438 9392 20444 9404
rect 20496 9432 20502 9444
rect 21266 9432 21272 9444
rect 20496 9404 21272 9432
rect 20496 9392 20502 9404
rect 21266 9392 21272 9404
rect 21324 9392 21330 9444
rect 17635 9336 18736 9364
rect 17635 9333 17647 9336
rect 17589 9327 17647 9333
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19521 9367 19579 9373
rect 19521 9364 19533 9367
rect 18932 9336 19533 9364
rect 18932 9324 18938 9336
rect 19521 9333 19533 9336
rect 19567 9333 19579 9367
rect 19521 9327 19579 9333
rect 21085 9367 21143 9373
rect 21085 9333 21097 9367
rect 21131 9364 21143 9367
rect 21174 9364 21180 9376
rect 21131 9336 21180 9364
rect 21131 9333 21143 9336
rect 21085 9327 21143 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21376 9364 21404 9540
rect 21450 9528 21456 9580
rect 21508 9528 21514 9580
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 22060 9540 22201 9568
rect 22060 9528 22066 9540
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9568 22339 9571
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22327 9540 22661 9568
rect 22327 9537 22339 9540
rect 22281 9531 22339 9537
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 22922 9528 22928 9580
rect 22980 9568 22986 9580
rect 23385 9571 23443 9577
rect 23385 9568 23397 9571
rect 22980 9540 23397 9568
rect 22980 9528 22986 9540
rect 23385 9537 23397 9540
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 21542 9460 21548 9512
rect 21600 9500 21606 9512
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 21600 9472 22385 9500
rect 21600 9460 21606 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 23201 9503 23259 9509
rect 23201 9469 23213 9503
rect 23247 9469 23259 9503
rect 23201 9463 23259 9469
rect 21637 9435 21695 9441
rect 21637 9401 21649 9435
rect 21683 9432 21695 9435
rect 21683 9404 22094 9432
rect 21683 9401 21695 9404
rect 21637 9395 21695 9401
rect 22066 9376 22094 9404
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 23216 9432 23244 9463
rect 22244 9404 23244 9432
rect 22244 9392 22250 9404
rect 23382 9392 23388 9444
rect 23440 9432 23446 9444
rect 23569 9435 23627 9441
rect 23569 9432 23581 9435
rect 23440 9404 23581 9432
rect 23440 9392 23446 9404
rect 23569 9401 23581 9404
rect 23615 9401 23627 9435
rect 23569 9395 23627 9401
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21376 9336 21833 9364
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 22066 9336 22100 9376
rect 21821 9327 21879 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 1104 9274 24012 9296
rect 1104 9222 1350 9274
rect 1402 9222 1414 9274
rect 1466 9222 1478 9274
rect 1530 9222 1542 9274
rect 1594 9222 1606 9274
rect 1658 9222 4350 9274
rect 4402 9222 4414 9274
rect 4466 9222 4478 9274
rect 4530 9222 4542 9274
rect 4594 9222 4606 9274
rect 4658 9222 7350 9274
rect 7402 9222 7414 9274
rect 7466 9222 7478 9274
rect 7530 9222 7542 9274
rect 7594 9222 7606 9274
rect 7658 9222 10350 9274
rect 10402 9222 10414 9274
rect 10466 9222 10478 9274
rect 10530 9222 10542 9274
rect 10594 9222 10606 9274
rect 10658 9222 13350 9274
rect 13402 9222 13414 9274
rect 13466 9222 13478 9274
rect 13530 9222 13542 9274
rect 13594 9222 13606 9274
rect 13658 9222 16350 9274
rect 16402 9222 16414 9274
rect 16466 9222 16478 9274
rect 16530 9222 16542 9274
rect 16594 9222 16606 9274
rect 16658 9222 19350 9274
rect 19402 9222 19414 9274
rect 19466 9222 19478 9274
rect 19530 9222 19542 9274
rect 19594 9222 19606 9274
rect 19658 9222 22350 9274
rect 22402 9222 22414 9274
rect 22466 9222 22478 9274
rect 22530 9222 22542 9274
rect 22594 9222 22606 9274
rect 22658 9222 24012 9274
rect 1104 9200 24012 9222
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 5810 9160 5816 9172
rect 5767 9132 5816 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 6454 9120 6460 9172
rect 6512 9120 6518 9172
rect 9674 9120 9680 9172
rect 9732 9120 9738 9172
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9129 10011 9163
rect 11514 9160 11520 9172
rect 9953 9123 10011 9129
rect 10244 9132 11520 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 3694 9092 3700 9104
rect 1627 9064 3004 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 382 8916 388 8968
rect 440 8956 446 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 440 8928 1409 8956
rect 440 8916 446 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8956 2467 8959
rect 2455 8928 2728 8956
rect 2455 8925 2467 8928
rect 2409 8919 2467 8925
rect 2222 8780 2228 8832
rect 2280 8780 2286 8832
rect 2700 8829 2728 8928
rect 2685 8823 2743 8829
rect 2685 8789 2697 8823
rect 2731 8789 2743 8823
rect 2976 8820 3004 9064
rect 3344 9064 3700 9092
rect 3344 9033 3372 9064
rect 3694 9052 3700 9064
rect 3752 9092 3758 9104
rect 5534 9092 5540 9104
rect 3752 9064 5540 9092
rect 3752 9052 3758 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 9769 9095 9827 9101
rect 9769 9092 9781 9095
rect 9416 9064 9781 9092
rect 9416 9036 9444 9064
rect 9769 9061 9781 9064
rect 9815 9061 9827 9095
rect 9769 9055 9827 9061
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 8993 3387 9027
rect 3329 8987 3387 8993
rect 5258 8984 5264 9036
rect 5316 8984 5322 9036
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5684 8996 6285 9024
rect 5684 8984 5690 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 7926 9024 7932 9036
rect 6273 8987 6331 8993
rect 6380 8996 7932 9024
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 3292 8928 4353 8956
rect 3292 8916 3298 8928
rect 4341 8925 4353 8928
rect 4387 8956 4399 8959
rect 4614 8956 4620 8968
rect 4387 8928 4620 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 5276 8956 5304 8984
rect 6380 8956 6408 8996
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9968 9024 9996 9123
rect 9640 8996 9996 9024
rect 9640 8984 9646 8996
rect 5276 8928 6408 8956
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 10244 8965 10272 9132
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 12434 9160 12440 9172
rect 12299 9132 12440 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12894 9160 12900 9172
rect 12544 9132 12900 9160
rect 10778 8984 10784 9036
rect 10836 8984 10842 9036
rect 12544 9033 12572 9132
rect 12894 9120 12900 9132
rect 12952 9160 12958 9172
rect 15194 9160 15200 9172
rect 12952 9132 15200 9160
rect 12952 9120 12958 9132
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 14108 9024 14136 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 15838 9160 15844 9172
rect 15611 9132 15844 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 18877 9163 18935 9169
rect 16264 9132 18460 9160
rect 16264 9120 16270 9132
rect 18432 9092 18460 9132
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19150 9160 19156 9172
rect 18923 9132 19156 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 19242 9120 19248 9172
rect 19300 9160 19306 9172
rect 20625 9163 20683 9169
rect 20625 9160 20637 9163
rect 19300 9132 20637 9160
rect 19300 9120 19306 9132
rect 20625 9129 20637 9132
rect 20671 9160 20683 9163
rect 20714 9160 20720 9172
rect 20671 9132 20720 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 22186 9120 22192 9172
rect 22244 9160 22250 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22244 9132 22293 9160
rect 22244 9120 22250 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 22833 9163 22891 9169
rect 22833 9129 22845 9163
rect 22879 9160 22891 9163
rect 22922 9160 22928 9172
rect 22879 9132 22928 9160
rect 22879 9129 22891 9132
rect 22833 9123 22891 9129
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 19058 9092 19064 9104
rect 18432 9064 19064 9092
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 22002 9052 22008 9104
rect 22060 9092 22066 9104
rect 23477 9095 23535 9101
rect 23477 9092 23489 9095
rect 22060 9064 23489 9092
rect 22060 9052 22066 9064
rect 23477 9061 23489 9064
rect 23523 9061 23535 9095
rect 23477 9055 23535 9061
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 14108 8996 14197 9024
rect 12529 8987 12587 8993
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 16022 9024 16028 9036
rect 15252 8996 16028 9024
rect 15252 8984 15258 8996
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 23290 8984 23296 9036
rect 23348 9024 23354 9036
rect 23348 8996 23704 9024
rect 23348 8984 23354 8996
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 8720 8928 9321 8956
rect 8720 8916 8726 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 3053 8891 3111 8897
rect 3053 8857 3065 8891
rect 3099 8888 3111 8891
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 3099 8860 3801 8888
rect 3099 8857 3111 8860
rect 3053 8851 3111 8857
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 3789 8851 3847 8857
rect 3988 8860 5028 8888
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 2976 8792 3157 8820
rect 2685 8783 2743 8789
rect 3145 8789 3157 8792
rect 3191 8820 3203 8823
rect 3988 8820 4016 8860
rect 5000 8832 5028 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 10520 8888 10548 8919
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 12785 8959 12843 8965
rect 12785 8956 12797 8959
rect 12676 8928 12797 8956
rect 12676 8916 12682 8928
rect 12785 8925 12797 8928
rect 12831 8925 12843 8959
rect 12785 8919 12843 8925
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 16908 8928 17509 8956
rect 16908 8916 16914 8928
rect 17497 8925 17509 8928
rect 17543 8956 17555 8959
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 17543 8928 19257 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 19245 8925 19257 8928
rect 19291 8956 19303 8959
rect 19794 8956 19800 8968
rect 19291 8928 19800 8956
rect 19291 8925 19303 8928
rect 19245 8919 19303 8925
rect 19794 8916 19800 8928
rect 19852 8956 19858 8968
rect 21174 8965 21180 8968
rect 20901 8959 20959 8965
rect 20901 8956 20913 8959
rect 19852 8928 20913 8956
rect 19852 8916 19858 8928
rect 20901 8925 20913 8928
rect 20947 8925 20959 8959
rect 21168 8956 21180 8965
rect 21135 8928 21180 8956
rect 20901 8919 20959 8925
rect 21168 8919 21180 8928
rect 21174 8916 21180 8919
rect 21232 8916 21238 8968
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8956 22707 8959
rect 22738 8956 22744 8968
rect 22695 8928 22744 8956
rect 22695 8925 22707 8928
rect 22649 8919 22707 8925
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 23382 8916 23388 8968
rect 23440 8916 23446 8968
rect 23676 8965 23704 8996
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 9548 8860 10548 8888
rect 9548 8848 9554 8860
rect 11514 8848 11520 8900
rect 11572 8848 11578 8900
rect 14452 8891 14510 8897
rect 14452 8857 14464 8891
rect 14498 8888 14510 8891
rect 14734 8888 14740 8900
rect 14498 8860 14740 8888
rect 14498 8857 14510 8860
rect 14452 8851 14510 8857
rect 14734 8848 14740 8860
rect 14792 8848 14798 8900
rect 16298 8897 16304 8900
rect 16292 8851 16304 8897
rect 16298 8848 16304 8851
rect 16356 8848 16362 8900
rect 17770 8897 17776 8900
rect 17764 8851 17776 8897
rect 17770 8848 17776 8851
rect 17828 8848 17834 8900
rect 18230 8848 18236 8900
rect 18288 8888 18294 8900
rect 19518 8897 19524 8900
rect 18288 8860 19334 8888
rect 18288 8848 18294 8860
rect 3191 8792 4016 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 4212 8792 4629 8820
rect 4212 8780 4218 8792
rect 4617 8789 4629 8792
rect 4663 8789 4675 8823
rect 4617 8783 4675 8789
rect 4982 8780 4988 8832
rect 5040 8780 5046 8832
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 6362 8820 6368 8832
rect 5123 8792 6368 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 8205 8823 8263 8829
rect 8205 8789 8217 8823
rect 8251 8820 8263 8823
rect 8294 8820 8300 8832
rect 8251 8792 8300 8820
rect 8251 8789 8263 8792
rect 8205 8783 8263 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 13909 8823 13967 8829
rect 13909 8789 13921 8823
rect 13955 8820 13967 8823
rect 14642 8820 14648 8832
rect 13955 8792 14648 8820
rect 13955 8789 13967 8792
rect 13909 8783 13967 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15841 8823 15899 8829
rect 15841 8789 15853 8823
rect 15887 8820 15899 8823
rect 16574 8820 16580 8832
rect 15887 8792 16580 8820
rect 15887 8789 15899 8792
rect 15841 8783 15899 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 18414 8820 18420 8832
rect 17451 8792 18420 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 19306 8820 19334 8860
rect 19512 8851 19524 8897
rect 19518 8848 19524 8851
rect 19576 8848 19582 8900
rect 21450 8888 21456 8900
rect 19628 8860 21456 8888
rect 19628 8820 19656 8860
rect 21450 8848 21456 8860
rect 21508 8848 21514 8900
rect 19306 8792 19656 8820
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 23201 8823 23259 8829
rect 23201 8820 23213 8823
rect 19944 8792 23213 8820
rect 19944 8780 19950 8792
rect 23201 8789 23213 8792
rect 23247 8789 23259 8823
rect 23201 8783 23259 8789
rect 1104 8730 24164 8752
rect 1104 8678 2850 8730
rect 2902 8678 2914 8730
rect 2966 8678 2978 8730
rect 3030 8678 3042 8730
rect 3094 8678 3106 8730
rect 3158 8678 5850 8730
rect 5902 8678 5914 8730
rect 5966 8678 5978 8730
rect 6030 8678 6042 8730
rect 6094 8678 6106 8730
rect 6158 8678 8850 8730
rect 8902 8678 8914 8730
rect 8966 8678 8978 8730
rect 9030 8678 9042 8730
rect 9094 8678 9106 8730
rect 9158 8678 11850 8730
rect 11902 8678 11914 8730
rect 11966 8678 11978 8730
rect 12030 8678 12042 8730
rect 12094 8678 12106 8730
rect 12158 8678 14850 8730
rect 14902 8678 14914 8730
rect 14966 8678 14978 8730
rect 15030 8678 15042 8730
rect 15094 8678 15106 8730
rect 15158 8678 17850 8730
rect 17902 8678 17914 8730
rect 17966 8678 17978 8730
rect 18030 8678 18042 8730
rect 18094 8678 18106 8730
rect 18158 8678 20850 8730
rect 20902 8678 20914 8730
rect 20966 8678 20978 8730
rect 21030 8678 21042 8730
rect 21094 8678 21106 8730
rect 21158 8678 23850 8730
rect 23902 8678 23914 8730
rect 23966 8678 23978 8730
rect 24030 8678 24042 8730
rect 24094 8678 24106 8730
rect 24158 8678 24164 8730
rect 1104 8656 24164 8678
rect 3234 8576 3240 8628
rect 3292 8576 3298 8628
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 3743 8588 5856 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 2124 8551 2182 8557
rect 2124 8517 2136 8551
rect 2170 8548 2182 8551
rect 2222 8548 2228 8560
rect 2170 8520 2228 8548
rect 2170 8517 2182 8520
rect 2124 8511 2182 8517
rect 2222 8508 2228 8520
rect 2280 8508 2286 8560
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1719 8452 3464 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 3436 8412 3464 8452
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4614 8440 4620 8492
rect 4672 8440 4678 8492
rect 5828 8489 5856 8588
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 9509 8619 9567 8625
rect 9509 8616 9521 8619
rect 9079 8588 9521 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9509 8585 9521 8588
rect 9555 8585 9567 8619
rect 9509 8579 9567 8585
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 10134 8616 10140 8628
rect 9723 8588 10140 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 13814 8576 13820 8628
rect 13872 8576 13878 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 14792 8588 15117 8616
rect 14792 8576 14798 8588
rect 15105 8585 15117 8588
rect 15151 8585 15163 8619
rect 15105 8579 15163 8585
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 16758 8576 16764 8628
rect 16816 8576 16822 8628
rect 17126 8576 17132 8628
rect 17184 8576 17190 8628
rect 17589 8619 17647 8625
rect 17589 8585 17601 8619
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 10042 8548 10048 8560
rect 9355 8520 10048 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 14921 8551 14979 8557
rect 14921 8517 14933 8551
rect 14967 8548 14979 8551
rect 15194 8548 15200 8560
rect 14967 8520 15200 8548
rect 14967 8517 14979 8520
rect 14921 8511 14979 8517
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 17604 8548 17632 8579
rect 18874 8576 18880 8628
rect 18932 8576 18938 8628
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 19518 8616 19524 8628
rect 19475 8588 19524 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 16500 8520 17632 8548
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5813 8483 5871 8489
rect 5399 8452 5764 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5736 8424 5764 8452
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 4522 8421 4528 8424
rect 4479 8415 4528 8421
rect 3436 8384 4016 8412
rect 1210 8304 1216 8356
rect 1268 8344 1274 8356
rect 1489 8347 1547 8353
rect 1489 8344 1501 8347
rect 1268 8316 1501 8344
rect 1268 8304 1274 8316
rect 1489 8313 1501 8316
rect 1535 8313 1547 8347
rect 1489 8307 1547 8313
rect 3326 8236 3332 8288
rect 3384 8236 3390 8288
rect 3988 8276 4016 8384
rect 4479 8381 4491 8415
rect 4525 8381 4528 8415
rect 4479 8375 4528 8381
rect 4522 8372 4528 8375
rect 4580 8372 4586 8424
rect 4890 8372 4896 8424
rect 4948 8372 4954 8424
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 5776 8384 6929 8412
rect 5776 8372 5782 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 4816 8316 5641 8344
rect 4816 8276 4844 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 8680 8344 8708 8443
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9272 8452 10149 8480
rect 9272 8440 9278 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 11698 8480 11704 8492
rect 10459 8452 11704 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 10336 8412 10364 8443
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14642 8480 14648 8492
rect 14507 8452 14648 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 16500 8489 16528 8520
rect 18046 8508 18052 8560
rect 18104 8508 18110 8560
rect 19705 8551 19763 8557
rect 19705 8517 19717 8551
rect 19751 8548 19763 8551
rect 19794 8548 19800 8560
rect 19751 8520 19800 8548
rect 19751 8517 19763 8520
rect 19705 8511 19763 8517
rect 19794 8508 19800 8520
rect 19852 8508 19858 8560
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17957 8483 18015 8489
rect 17957 8480 17969 8483
rect 17267 8452 17969 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17957 8449 17969 8452
rect 18003 8480 18015 8483
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18003 8452 18797 8480
rect 18003 8449 18015 8452
rect 17957 8443 18015 8449
rect 18785 8449 18797 8452
rect 18831 8480 18843 8483
rect 18831 8452 19196 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 9364 8384 10364 8412
rect 9364 8372 9370 8384
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 14608 8384 17325 8412
rect 14608 8372 14614 8384
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17920 8384 18153 8412
rect 17920 8372 17926 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 19061 8415 19119 8421
rect 19061 8381 19073 8415
rect 19107 8381 19119 8415
rect 19168 8412 19196 8452
rect 19242 8440 19248 8492
rect 19300 8440 19306 8492
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8480 20499 8483
rect 20622 8480 20628 8492
rect 20487 8452 20628 8480
rect 20487 8449 20499 8452
rect 20441 8443 20499 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 21085 8483 21143 8489
rect 21085 8480 21097 8483
rect 20772 8452 21097 8480
rect 20772 8440 20778 8452
rect 21085 8449 21097 8452
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 19886 8412 19892 8424
rect 19168 8384 19892 8412
rect 19061 8375 19119 8381
rect 5629 8307 5687 8313
rect 5736 8316 8708 8344
rect 3988 8248 4844 8276
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5736 8276 5764 8316
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 19076 8344 19104 8375
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 20714 8344 20720 8356
rect 16632 8316 20720 8344
rect 16632 8304 16638 8316
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 4948 8248 5764 8276
rect 4948 8236 4954 8248
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 6972 8248 7849 8276
rect 6972 8236 6978 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 7837 8239 7895 8245
rect 9398 8236 9404 8288
rect 9456 8276 9462 8288
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 9456 8248 9505 8276
rect 9456 8236 9462 8248
rect 9493 8245 9505 8248
rect 9539 8245 9551 8279
rect 9493 8239 9551 8245
rect 10134 8236 10140 8288
rect 10192 8236 10198 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18417 8279 18475 8285
rect 18417 8276 18429 8279
rect 18012 8248 18429 8276
rect 18012 8236 18018 8248
rect 18417 8245 18429 8248
rect 18463 8245 18475 8279
rect 18417 8239 18475 8245
rect 19702 8236 19708 8288
rect 19760 8276 19766 8288
rect 20533 8279 20591 8285
rect 20533 8276 20545 8279
rect 19760 8248 20545 8276
rect 19760 8236 19766 8248
rect 20533 8245 20545 8248
rect 20579 8245 20591 8279
rect 20533 8239 20591 8245
rect 1104 8186 24012 8208
rect 1104 8134 1350 8186
rect 1402 8134 1414 8186
rect 1466 8134 1478 8186
rect 1530 8134 1542 8186
rect 1594 8134 1606 8186
rect 1658 8134 4350 8186
rect 4402 8134 4414 8186
rect 4466 8134 4478 8186
rect 4530 8134 4542 8186
rect 4594 8134 4606 8186
rect 4658 8134 7350 8186
rect 7402 8134 7414 8186
rect 7466 8134 7478 8186
rect 7530 8134 7542 8186
rect 7594 8134 7606 8186
rect 7658 8134 10350 8186
rect 10402 8134 10414 8186
rect 10466 8134 10478 8186
rect 10530 8134 10542 8186
rect 10594 8134 10606 8186
rect 10658 8134 13350 8186
rect 13402 8134 13414 8186
rect 13466 8134 13478 8186
rect 13530 8134 13542 8186
rect 13594 8134 13606 8186
rect 13658 8134 16350 8186
rect 16402 8134 16414 8186
rect 16466 8134 16478 8186
rect 16530 8134 16542 8186
rect 16594 8134 16606 8186
rect 16658 8134 19350 8186
rect 19402 8134 19414 8186
rect 19466 8134 19478 8186
rect 19530 8134 19542 8186
rect 19594 8134 19606 8186
rect 19658 8134 22350 8186
rect 22402 8134 22414 8186
rect 22466 8134 22478 8186
rect 22530 8134 22542 8186
rect 22594 8134 22606 8186
rect 22658 8134 24012 8186
rect 1104 8112 24012 8134
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 3844 8044 5825 8072
rect 3844 8032 3850 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 8076 8044 8125 8072
rect 8076 8032 8082 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 9214 8072 9220 8084
rect 8343 8044 9220 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 3237 8007 3295 8013
rect 3237 7973 3249 8007
rect 3283 8004 3295 8007
rect 4338 8004 4344 8016
rect 3283 7976 4344 8004
rect 3283 7973 3295 7976
rect 3237 7967 3295 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 5718 7964 5724 8016
rect 5776 7964 5782 8016
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8312 8004 8340 8035
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 13081 8075 13139 8081
rect 13081 8041 13093 8075
rect 13127 8072 13139 8075
rect 13262 8072 13268 8084
rect 13127 8044 13268 8072
rect 13127 8041 13139 8044
rect 13081 8035 13139 8041
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 17770 8072 17776 8084
rect 17727 8044 17776 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 19242 8032 19248 8084
rect 19300 8032 19306 8084
rect 20714 8072 20720 8084
rect 20180 8044 20720 8072
rect 7984 7976 8340 8004
rect 7984 7964 7990 7976
rect 10134 7964 10140 8016
rect 10192 7964 10198 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 14645 8007 14703 8013
rect 12676 7976 13676 8004
rect 12676 7964 12682 7976
rect 6457 7939 6515 7945
rect 3712 7908 4384 7936
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 3712 7868 3740 7908
rect 4356 7880 4384 7908
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 8110 7936 8116 7948
rect 6503 7908 7512 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 1912 7840 3740 7868
rect 1912 7828 1918 7840
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4154 7868 4160 7880
rect 4111 7840 4160 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 5534 7828 5540 7880
rect 5592 7868 5598 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 5592 7840 7205 7868
rect 5592 7828 5598 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 2124 7803 2182 7809
rect 2124 7769 2136 7803
rect 2170 7800 2182 7803
rect 3326 7800 3332 7812
rect 2170 7772 3332 7800
rect 2170 7769 2182 7772
rect 2124 7763 2182 7769
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 4586 7803 4644 7809
rect 4586 7800 4598 7803
rect 4264 7772 4598 7800
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 4264 7741 4292 7772
rect 4586 7769 4598 7772
rect 4632 7769 4644 7803
rect 4586 7763 4644 7769
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 6181 7803 6239 7809
rect 6181 7800 6193 7803
rect 5040 7772 6193 7800
rect 5040 7760 5046 7772
rect 6181 7769 6193 7772
rect 6227 7769 6239 7803
rect 6181 7763 6239 7769
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 6319 7704 6653 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6641 7701 6653 7704
rect 6687 7701 6699 7735
rect 6641 7695 6699 7701
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 6972 7704 7389 7732
rect 6972 7692 6978 7704
rect 7377 7701 7389 7704
rect 7423 7701 7435 7735
rect 7484 7732 7512 7908
rect 7668 7908 8116 7936
rect 7668 7877 7696 7908
rect 8110 7896 8116 7908
rect 8168 7936 8174 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8168 7908 8401 7936
rect 8168 7896 8174 7908
rect 8389 7905 8401 7908
rect 8435 7936 8447 7939
rect 8846 7936 8852 7948
rect 8435 7908 8852 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 10152 7936 10180 7964
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 10152 7908 10425 7936
rect 10413 7905 10425 7908
rect 10459 7905 10471 7939
rect 10413 7899 10471 7905
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12529 7939 12587 7945
rect 12529 7936 12541 7939
rect 11931 7908 12541 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12529 7905 12541 7908
rect 12575 7936 12587 7939
rect 12575 7908 12940 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7576 7800 7604 7831
rect 7742 7800 7748 7812
rect 7576 7772 7748 7800
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 7852 7800 7880 7831
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 9214 7868 9220 7880
rect 8711 7840 9220 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9548 7840 10149 7868
rect 9548 7828 9554 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 12912 7877 12940 7908
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 13170 7868 13176 7880
rect 12943 7840 13176 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13648 7877 13676 7976
rect 14645 7973 14657 8007
rect 14691 8004 14703 8007
rect 17218 8004 17224 8016
rect 14691 7976 17224 8004
rect 14691 7973 14703 7976
rect 14645 7967 14703 7973
rect 17218 7964 17224 7976
rect 17276 8004 17282 8016
rect 17276 7976 19840 8004
rect 17276 7964 17282 7976
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7936 17831 7939
rect 18046 7936 18052 7948
rect 17819 7908 18052 7936
rect 17819 7905 17831 7908
rect 17773 7899 17831 7905
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18414 7896 18420 7948
rect 18472 7896 18478 7948
rect 19702 7896 19708 7948
rect 19760 7896 19766 7948
rect 19812 7945 19840 7976
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 20180 7936 20208 8044
rect 20714 8032 20720 8044
rect 20772 8072 20778 8084
rect 21542 8072 21548 8084
rect 20772 8044 21548 8072
rect 20772 8032 20778 8044
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 20257 8007 20315 8013
rect 20257 7973 20269 8007
rect 20303 8004 20315 8007
rect 21818 8004 21824 8016
rect 20303 7976 21824 8004
rect 20303 7973 20315 7976
rect 20257 7967 20315 7973
rect 21818 7964 21824 7976
rect 21876 7964 21882 8016
rect 20441 7939 20499 7945
rect 20441 7936 20453 7939
rect 20036 7908 20453 7936
rect 20036 7896 20042 7908
rect 20441 7905 20453 7908
rect 20487 7905 20499 7939
rect 20441 7899 20499 7905
rect 20530 7896 20536 7948
rect 20588 7936 20594 7948
rect 21729 7939 21787 7945
rect 21729 7936 21741 7939
rect 20588 7908 21741 7936
rect 20588 7896 20594 7908
rect 21729 7905 21741 7908
rect 21775 7905 21787 7939
rect 21729 7899 21787 7905
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14274 7828 14280 7880
rect 14332 7868 14338 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14332 7840 14473 7868
rect 14332 7828 14338 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7868 17555 7871
rect 17954 7868 17960 7880
rect 17543 7840 17960 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 19886 7868 19892 7880
rect 19659 7840 19892 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7868 20131 7871
rect 21266 7868 21272 7880
rect 20119 7840 21272 7868
rect 20119 7837 20131 7840
rect 20073 7831 20131 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 8202 7800 8208 7812
rect 7852 7772 8208 7800
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 12710 7760 12716 7812
rect 12768 7760 12774 7812
rect 20625 7803 20683 7809
rect 20625 7769 20637 7803
rect 20671 7800 20683 7803
rect 21177 7803 21235 7809
rect 21177 7800 21189 7803
rect 20671 7772 21189 7800
rect 20671 7769 20683 7772
rect 20625 7763 20683 7769
rect 21177 7769 21189 7772
rect 21223 7769 21235 7803
rect 21177 7763 21235 7769
rect 9306 7732 9312 7744
rect 7484 7704 9312 7732
rect 7377 7695 7435 7701
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12250 7732 12256 7744
rect 12023 7704 12256 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 13814 7692 13820 7744
rect 13872 7692 13878 7744
rect 14277 7735 14335 7741
rect 14277 7701 14289 7735
rect 14323 7732 14335 7735
rect 14550 7732 14556 7744
rect 14323 7704 14556 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 20714 7692 20720 7744
rect 20772 7692 20778 7744
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 1104 7642 24164 7664
rect 1104 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 3042 7642
rect 3094 7590 3106 7642
rect 3158 7590 5850 7642
rect 5902 7590 5914 7642
rect 5966 7590 5978 7642
rect 6030 7590 6042 7642
rect 6094 7590 6106 7642
rect 6158 7590 8850 7642
rect 8902 7590 8914 7642
rect 8966 7590 8978 7642
rect 9030 7590 9042 7642
rect 9094 7590 9106 7642
rect 9158 7590 11850 7642
rect 11902 7590 11914 7642
rect 11966 7590 11978 7642
rect 12030 7590 12042 7642
rect 12094 7590 12106 7642
rect 12158 7590 14850 7642
rect 14902 7590 14914 7642
rect 14966 7590 14978 7642
rect 15030 7590 15042 7642
rect 15094 7590 15106 7642
rect 15158 7590 17850 7642
rect 17902 7590 17914 7642
rect 17966 7590 17978 7642
rect 18030 7590 18042 7642
rect 18094 7590 18106 7642
rect 18158 7590 20850 7642
rect 20902 7590 20914 7642
rect 20966 7590 20978 7642
rect 21030 7590 21042 7642
rect 21094 7590 21106 7642
rect 21158 7590 23850 7642
rect 23902 7590 23914 7642
rect 23966 7590 23978 7642
rect 24030 7590 24042 7642
rect 24094 7590 24106 7642
rect 24158 7590 24164 7642
rect 1104 7568 24164 7590
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3510 7528 3516 7540
rect 3375 7500 3516 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5534 7528 5540 7540
rect 5399 7500 5540 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 8260 7500 8401 7528
rect 8260 7488 8266 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 8389 7491 8447 7497
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 11756 7500 12081 7528
rect 11756 7488 11762 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 14274 7528 14280 7540
rect 13679 7500 14280 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 19852 7500 20269 7528
rect 19852 7488 19858 7500
rect 20257 7497 20269 7500
rect 20303 7528 20315 7531
rect 20530 7528 20536 7540
rect 20303 7500 20536 7528
rect 20303 7497 20315 7500
rect 20257 7491 20315 7497
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21542 7528 21548 7540
rect 20772 7500 21548 7528
rect 20772 7488 20778 7500
rect 21542 7488 21548 7500
rect 21600 7488 21606 7540
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4218 7463 4276 7469
rect 4218 7460 4230 7463
rect 4028 7432 4230 7460
rect 4028 7420 4034 7432
rect 4218 7429 4230 7432
rect 4264 7429 4276 7463
rect 4218 7423 4276 7429
rect 7190 7420 7196 7472
rect 7248 7420 7254 7472
rect 12710 7460 12716 7472
rect 8404 7432 8800 7460
rect 8404 7404 8432 7432
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 4982 7392 4988 7404
rect 3007 7364 4988 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 6472 7364 6960 7392
rect 2774 7284 2780 7336
rect 2832 7284 2838 7336
rect 2866 7284 2872 7336
rect 2924 7284 2930 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 3988 7188 4016 7287
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 6472 7333 6500 7364
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 6236 7296 6469 7324
rect 6236 7284 6242 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 6932 7324 6960 7364
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8772 7401 8800 7432
rect 9048 7432 9352 7460
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8536 7364 8677 7392
rect 8536 7352 8542 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 9048 7401 9076 7432
rect 9324 7404 9352 7432
rect 11992 7432 12716 7460
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9214 7392 9220 7404
rect 9171 7364 9220 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9582 7392 9588 7404
rect 9364 7364 9588 7392
rect 9364 7352 9370 7364
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 11992 7401 12020 7432
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 15194 7420 15200 7472
rect 15252 7420 15258 7472
rect 19153 7463 19211 7469
rect 19153 7429 19165 7463
rect 19199 7460 19211 7463
rect 21821 7463 21879 7469
rect 21821 7460 21833 7463
rect 19199 7432 21833 7460
rect 19199 7429 19211 7432
rect 19153 7423 19211 7429
rect 21821 7429 21833 7432
rect 21867 7429 21879 7463
rect 21821 7423 21879 7429
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12250 7392 12256 7404
rect 12207 7364 12256 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12805 7395 12863 7401
rect 12805 7392 12817 7395
rect 12492 7364 12817 7392
rect 12492 7352 12498 7364
rect 12805 7361 12817 7364
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 8294 7324 8300 7336
rect 6932 7296 8300 7324
rect 8294 7284 8300 7296
rect 8352 7324 8358 7336
rect 9490 7324 9496 7336
rect 8352 7296 9496 7324
rect 8352 7284 8358 7296
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 12820 7324 12848 7355
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 13228 7364 13277 7392
rect 13228 7352 13234 7364
rect 13265 7361 13277 7364
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 16850 7352 16856 7404
rect 16908 7392 16914 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16908 7364 17049 7392
rect 16908 7352 16914 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 17175 7364 17509 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 17678 7352 17684 7404
rect 17736 7392 17742 7404
rect 18417 7395 18475 7401
rect 18417 7392 18429 7395
rect 17736 7364 18429 7392
rect 17736 7352 17742 7364
rect 18417 7361 18429 7364
rect 18463 7361 18475 7395
rect 18417 7355 18475 7361
rect 19058 7352 19064 7404
rect 19116 7392 19122 7404
rect 20806 7392 20812 7404
rect 19116 7364 20812 7392
rect 19116 7352 19122 7364
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 21358 7352 21364 7404
rect 21416 7401 21422 7404
rect 21416 7355 21428 7401
rect 21416 7352 21422 7355
rect 22830 7352 22836 7404
rect 22888 7392 22894 7404
rect 23385 7395 23443 7401
rect 23385 7392 23397 7395
rect 22888 7364 23397 7392
rect 22888 7352 22894 7364
rect 23385 7361 23397 7364
rect 23431 7361 23443 7395
rect 23385 7355 23443 7361
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 12820 7296 13369 7324
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7324 13967 7327
rect 14458 7324 14464 7336
rect 13955 7296 14464 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15470 7284 15476 7336
rect 15528 7324 15534 7336
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 15528 7296 16313 7324
rect 15528 7284 15534 7296
rect 16301 7293 16313 7296
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 18012 7296 18061 7324
rect 18012 7284 18018 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 19245 7327 19303 7333
rect 19245 7293 19257 7327
rect 19291 7293 19303 7327
rect 19245 7287 19303 7293
rect 15562 7216 15568 7268
rect 15620 7256 15626 7268
rect 17770 7256 17776 7268
rect 15620 7228 17776 7256
rect 15620 7216 15626 7228
rect 17770 7216 17776 7228
rect 17828 7256 17834 7268
rect 19260 7256 19288 7287
rect 20070 7284 20076 7336
rect 20128 7284 20134 7336
rect 21634 7284 21640 7336
rect 21692 7284 21698 7336
rect 21726 7284 21732 7336
rect 21784 7324 21790 7336
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 21784 7296 22385 7324
rect 21784 7284 21790 7296
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 17828 7228 19288 7256
rect 17828 7216 17834 7228
rect 4338 7188 4344 7200
rect 3988 7160 4344 7188
rect 4338 7148 4344 7160
rect 4396 7188 4402 7200
rect 4706 7188 4712 7200
rect 4396 7160 4712 7188
rect 4396 7148 4402 7160
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 8251 7191 8309 7197
rect 8251 7157 8263 7191
rect 8297 7188 8309 7191
rect 8570 7188 8576 7200
rect 8297 7160 8576 7188
rect 8297 7157 8309 7160
rect 8251 7151 8309 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 9122 7148 9128 7200
rect 9180 7148 9186 7200
rect 13081 7191 13139 7197
rect 13081 7157 13093 7191
rect 13127 7188 13139 7191
rect 13262 7188 13268 7200
rect 13127 7160 13268 7188
rect 13127 7157 13139 7160
rect 13081 7151 13139 7157
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 15746 7148 15752 7200
rect 15804 7148 15810 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 16172 7160 16681 7188
rect 16172 7148 16178 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 18233 7191 18291 7197
rect 18233 7157 18245 7191
rect 18279 7188 18291 7191
rect 18414 7188 18420 7200
rect 18279 7160 18420 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18693 7191 18751 7197
rect 18693 7157 18705 7191
rect 18739 7188 18751 7191
rect 18782 7188 18788 7200
rect 18739 7160 18788 7188
rect 18739 7157 18751 7160
rect 18693 7151 18751 7157
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 19521 7191 19579 7197
rect 19521 7157 19533 7191
rect 19567 7188 19579 7191
rect 19702 7188 19708 7200
rect 19567 7160 19708 7188
rect 19567 7157 19579 7160
rect 19521 7151 19579 7157
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 23382 7148 23388 7200
rect 23440 7188 23446 7200
rect 23569 7191 23627 7197
rect 23569 7188 23581 7191
rect 23440 7160 23581 7188
rect 23440 7148 23446 7160
rect 23569 7157 23581 7160
rect 23615 7157 23627 7191
rect 23569 7151 23627 7157
rect 1104 7098 24012 7120
rect 1104 7046 1350 7098
rect 1402 7046 1414 7098
rect 1466 7046 1478 7098
rect 1530 7046 1542 7098
rect 1594 7046 1606 7098
rect 1658 7046 4350 7098
rect 4402 7046 4414 7098
rect 4466 7046 4478 7098
rect 4530 7046 4542 7098
rect 4594 7046 4606 7098
rect 4658 7046 7350 7098
rect 7402 7046 7414 7098
rect 7466 7046 7478 7098
rect 7530 7046 7542 7098
rect 7594 7046 7606 7098
rect 7658 7046 10350 7098
rect 10402 7046 10414 7098
rect 10466 7046 10478 7098
rect 10530 7046 10542 7098
rect 10594 7046 10606 7098
rect 10658 7046 13350 7098
rect 13402 7046 13414 7098
rect 13466 7046 13478 7098
rect 13530 7046 13542 7098
rect 13594 7046 13606 7098
rect 13658 7046 16350 7098
rect 16402 7046 16414 7098
rect 16466 7046 16478 7098
rect 16530 7046 16542 7098
rect 16594 7046 16606 7098
rect 16658 7046 19350 7098
rect 19402 7046 19414 7098
rect 19466 7046 19478 7098
rect 19530 7046 19542 7098
rect 19594 7046 19606 7098
rect 19658 7046 22350 7098
rect 22402 7046 22414 7098
rect 22466 7046 22478 7098
rect 22530 7046 22542 7098
rect 22594 7046 22606 7098
rect 22658 7046 24012 7098
rect 1104 7024 24012 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 2924 6956 3801 6984
rect 2924 6944 2930 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 3789 6947 3847 6953
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8021 6987 8079 6993
rect 8021 6984 8033 6987
rect 7800 6956 8033 6984
rect 7800 6944 7806 6956
rect 8021 6953 8033 6956
rect 8067 6953 8079 6987
rect 8021 6947 8079 6953
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9493 6987 9551 6993
rect 9493 6984 9505 6987
rect 9180 6956 9505 6984
rect 9180 6944 9186 6956
rect 9493 6953 9505 6956
rect 9539 6953 9551 6987
rect 9493 6947 9551 6953
rect 11793 6987 11851 6993
rect 11793 6953 11805 6987
rect 11839 6984 11851 6987
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 11839 6956 12265 6984
rect 11839 6953 11851 6956
rect 11793 6947 11851 6953
rect 12253 6953 12265 6956
rect 12299 6984 12311 6987
rect 12710 6984 12716 6996
rect 12299 6956 12716 6984
rect 12299 6953 12311 6956
rect 12253 6947 12311 6953
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 12897 6987 12955 6993
rect 12897 6953 12909 6987
rect 12943 6984 12955 6987
rect 13262 6984 13268 6996
rect 12943 6956 13268 6984
rect 12943 6953 12955 6956
rect 12897 6947 12955 6953
rect 7834 6876 7840 6928
rect 7892 6916 7898 6928
rect 7892 6888 9628 6916
rect 7892 6876 7898 6888
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 4304 6820 4353 6848
rect 4304 6808 4310 6820
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 6914 6848 6920 6860
rect 6503 6820 6920 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 9600 6857 9628 6888
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8720 6820 9045 6848
rect 8720 6808 8726 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 9033 6811 9091 6817
rect 9140 6820 9229 6848
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6178 6780 6184 6792
rect 6135 6752 6184 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8496 6752 8953 6780
rect 7190 6672 7196 6724
rect 7248 6672 7254 6724
rect 7883 6647 7941 6653
rect 7883 6613 7895 6647
rect 7929 6644 7941 6647
rect 8018 6644 8024 6656
rect 7929 6616 8024 6644
rect 7929 6613 7941 6616
rect 7883 6607 7941 6613
rect 8018 6604 8024 6616
rect 8076 6644 8082 6656
rect 8386 6644 8392 6656
rect 8076 6616 8392 6644
rect 8076 6604 8082 6616
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8496 6653 8524 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 8570 6672 8576 6724
rect 8628 6712 8634 6724
rect 9140 6712 9168 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 9631 6820 10149 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 12912 6848 12940 6947
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 21726 6984 21732 6996
rect 20956 6956 21732 6984
rect 20956 6944 20962 6956
rect 21726 6944 21732 6956
rect 21784 6944 21790 6996
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 15562 6916 15568 6928
rect 13872 6888 15568 6916
rect 13872 6876 13878 6888
rect 15212 6857 15240 6888
rect 15562 6876 15568 6888
rect 15620 6876 15626 6928
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 20128 6888 20576 6916
rect 20128 6876 20134 6888
rect 10137 6811 10195 6817
rect 10244 6820 11744 6848
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 8628 6684 9168 6712
rect 8628 6672 8634 6684
rect 9214 6672 9220 6724
rect 9272 6672 9278 6724
rect 9508 6712 9536 6743
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10244 6780 10272 6820
rect 11716 6792 11744 6820
rect 12360 6820 12940 6848
rect 15197 6851 15255 6857
rect 10100 6752 10272 6780
rect 11333 6783 11391 6789
rect 10100 6740 10106 6752
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11379 6752 11652 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 9766 6712 9772 6724
rect 9508 6684 9772 6712
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 9674 6644 9680 6656
rect 8527 6616 9680 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 10042 6644 10048 6656
rect 9907 6616 10048 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 11514 6604 11520 6656
rect 11572 6604 11578 6656
rect 11624 6653 11652 6752
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 12360 6789 12388 6820
rect 15197 6817 15209 6851
rect 15243 6817 15255 6851
rect 15654 6848 15660 6860
rect 15197 6811 15255 6817
rect 15304 6820 15660 6848
rect 12344 6783 12402 6789
rect 12344 6749 12356 6783
rect 12390 6749 12402 6783
rect 12344 6743 12402 6749
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 15304 6780 15332 6820
rect 15654 6808 15660 6820
rect 15712 6848 15718 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15712 6820 16037 6848
rect 15712 6808 15718 6820
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16025 6811 16083 6817
rect 18874 6808 18880 6860
rect 18932 6808 18938 6860
rect 19702 6808 19708 6860
rect 19760 6808 19766 6860
rect 19794 6808 19800 6860
rect 19852 6808 19858 6860
rect 20438 6808 20444 6860
rect 20496 6808 20502 6860
rect 20548 6848 20576 6888
rect 21450 6876 21456 6928
rect 21508 6876 21514 6928
rect 20898 6857 20904 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 20548 6820 20729 6848
rect 20717 6817 20729 6820
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20855 6851 20904 6857
rect 20855 6817 20867 6851
rect 20901 6817 20904 6851
rect 20855 6811 20904 6817
rect 20898 6808 20904 6811
rect 20956 6808 20962 6860
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 21468 6848 21496 6876
rect 21039 6820 21496 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 14516 6752 15332 6780
rect 15749 6783 15807 6789
rect 14516 6740 14522 6752
rect 15749 6749 15761 6783
rect 15795 6780 15807 6783
rect 16758 6780 16764 6792
rect 15795 6752 16764 6780
rect 15795 6749 15807 6752
rect 15749 6743 15807 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17644 6752 18061 6780
rect 17644 6740 17650 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 19720 6780 19748 6808
rect 18739 6752 19748 6780
rect 19981 6783 20039 6789
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 19981 6749 19993 6783
rect 20027 6780 20039 6783
rect 20162 6780 20168 6792
rect 20027 6752 20168 6780
rect 20027 6749 20039 6752
rect 19981 6743 20039 6749
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 21634 6780 21640 6792
rect 21560 6752 21640 6780
rect 11716 6712 11744 6740
rect 11977 6715 12035 6721
rect 11977 6712 11989 6715
rect 11716 6684 11989 6712
rect 11977 6681 11989 6684
rect 12023 6681 12035 6715
rect 11977 6675 12035 6681
rect 12526 6672 12532 6724
rect 12584 6712 12590 6724
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 12584 6684 12725 6712
rect 12584 6672 12590 6684
rect 12713 6681 12725 6684
rect 12759 6681 12771 6715
rect 12713 6675 12771 6681
rect 12929 6715 12987 6721
rect 12929 6681 12941 6715
rect 12975 6712 12987 6715
rect 13170 6712 13176 6724
rect 12975 6684 13176 6712
rect 12975 6681 12987 6684
rect 12929 6675 12987 6681
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 13998 6712 14004 6724
rect 13648 6684 14004 6712
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6613 11667 6647
rect 11609 6607 11667 6613
rect 11777 6647 11835 6653
rect 11777 6613 11789 6647
rect 11823 6644 11835 6647
rect 12342 6644 12348 6656
rect 11823 6616 12348 6644
rect 11823 6613 11835 6616
rect 11777 6607 11835 6613
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 13081 6647 13139 6653
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13648 6644 13676 6684
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 15013 6715 15071 6721
rect 15013 6681 15025 6715
rect 15059 6712 15071 6715
rect 15194 6712 15200 6724
rect 15059 6684 15200 6712
rect 15059 6681 15071 6684
rect 15013 6675 15071 6681
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 16292 6715 16350 6721
rect 16292 6681 16304 6715
rect 16338 6681 16350 6715
rect 17954 6712 17960 6724
rect 16292 6675 16350 6681
rect 17420 6684 17960 6712
rect 13127 6616 13676 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 13872 6616 14657 6644
rect 13872 6604 13878 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 15105 6647 15163 6653
rect 15105 6613 15117 6647
rect 15151 6644 15163 6647
rect 15286 6644 15292 6656
rect 15151 6616 15292 6644
rect 15151 6613 15163 6616
rect 15105 6607 15163 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16022 6644 16028 6656
rect 15979 6616 16028 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 16316 6644 16344 6675
rect 17420 6653 17448 6684
rect 17954 6672 17960 6684
rect 18012 6712 18018 6724
rect 18230 6712 18236 6724
rect 18012 6684 18236 6712
rect 18012 6672 18018 6684
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 18785 6715 18843 6721
rect 18785 6681 18797 6715
rect 18831 6712 18843 6715
rect 19058 6712 19064 6724
rect 18831 6684 19064 6712
rect 18831 6681 18843 6684
rect 18785 6675 18843 6681
rect 19058 6672 19064 6684
rect 19116 6672 19122 6724
rect 19337 6715 19395 6721
rect 19337 6681 19349 6715
rect 19383 6712 19395 6715
rect 19702 6712 19708 6724
rect 19383 6684 19708 6712
rect 19383 6681 19395 6684
rect 19337 6675 19395 6681
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 16264 6616 16344 6644
rect 17405 6647 17463 6653
rect 16264 6604 16270 6616
rect 17405 6613 17417 6647
rect 17451 6613 17463 6647
rect 17405 6607 17463 6613
rect 17494 6604 17500 6656
rect 17552 6604 17558 6656
rect 18322 6604 18328 6656
rect 18380 6604 18386 6656
rect 19720 6644 19748 6672
rect 21560 6644 21588 6752
rect 21634 6740 21640 6752
rect 21692 6780 21698 6792
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21692 6752 21741 6780
rect 21692 6740 21698 6752
rect 21729 6749 21741 6752
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 21818 6740 21824 6792
rect 21876 6780 21882 6792
rect 21985 6783 22043 6789
rect 21985 6780 21997 6783
rect 21876 6752 21997 6780
rect 21876 6740 21882 6752
rect 21985 6749 21997 6752
rect 22031 6749 22043 6783
rect 21985 6743 22043 6749
rect 19720 6616 21588 6644
rect 21634 6604 21640 6656
rect 21692 6604 21698 6656
rect 23106 6604 23112 6656
rect 23164 6604 23170 6656
rect 1104 6554 24164 6576
rect 1104 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 3042 6554
rect 3094 6502 3106 6554
rect 3158 6502 5850 6554
rect 5902 6502 5914 6554
rect 5966 6502 5978 6554
rect 6030 6502 6042 6554
rect 6094 6502 6106 6554
rect 6158 6502 8850 6554
rect 8902 6502 8914 6554
rect 8966 6502 8978 6554
rect 9030 6502 9042 6554
rect 9094 6502 9106 6554
rect 9158 6502 11850 6554
rect 11902 6502 11914 6554
rect 11966 6502 11978 6554
rect 12030 6502 12042 6554
rect 12094 6502 12106 6554
rect 12158 6502 14850 6554
rect 14902 6502 14914 6554
rect 14966 6502 14978 6554
rect 15030 6502 15042 6554
rect 15094 6502 15106 6554
rect 15158 6502 17850 6554
rect 17902 6502 17914 6554
rect 17966 6502 17978 6554
rect 18030 6502 18042 6554
rect 18094 6502 18106 6554
rect 18158 6502 20850 6554
rect 20902 6502 20914 6554
rect 20966 6502 20978 6554
rect 21030 6502 21042 6554
rect 21094 6502 21106 6554
rect 21158 6502 23850 6554
rect 23902 6502 23914 6554
rect 23966 6502 23978 6554
rect 24030 6502 24042 6554
rect 24094 6502 24106 6554
rect 24158 6502 24164 6554
rect 1104 6480 24164 6502
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 8168 6412 8217 6440
rect 8168 6400 8174 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 8205 6403 8263 6409
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 11054 6440 11060 6452
rect 10192 6412 11060 6440
rect 10192 6400 10198 6412
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 11606 6440 11612 6452
rect 11348 6412 11612 6440
rect 11348 6372 11376 6412
rect 11606 6400 11612 6412
rect 11664 6440 11670 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 11664 6412 11928 6440
rect 11664 6400 11670 6412
rect 10902 6344 11376 6372
rect 11514 6332 11520 6384
rect 11572 6372 11578 6384
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11572 6344 11805 6372
rect 11572 6332 11578 6344
rect 11793 6341 11805 6344
rect 11839 6341 11851 6375
rect 11900 6372 11928 6412
rect 13556 6412 15577 6440
rect 12250 6372 12256 6384
rect 11900 6344 12256 6372
rect 11793 6335 11851 6341
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 9122 6304 9128 6316
rect 8711 6276 9128 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 8312 6236 8340 6267
rect 9122 6264 9128 6276
rect 9180 6304 9186 6316
rect 9306 6304 9312 6316
rect 9180 6276 9312 6304
rect 9180 6264 9186 6276
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 13556 6313 13584 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15804 6412 15945 6440
rect 15804 6400 15810 6412
rect 15933 6409 15945 6412
rect 15979 6409 15991 6443
rect 15933 6403 15991 6409
rect 16669 6443 16727 6449
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 17586 6440 17592 6452
rect 16715 6412 17592 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 19613 6443 19671 6449
rect 19613 6409 19625 6443
rect 19659 6440 19671 6443
rect 20070 6440 20076 6452
rect 19659 6412 20076 6440
rect 19659 6409 19671 6412
rect 19613 6403 19671 6409
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 21358 6400 21364 6452
rect 21416 6400 21422 6452
rect 21637 6443 21695 6449
rect 21637 6409 21649 6443
rect 21683 6440 21695 6443
rect 22830 6440 22836 6452
rect 21683 6412 22836 6440
rect 21683 6409 21695 6412
rect 21637 6403 21695 6409
rect 22830 6400 22836 6412
rect 22888 6400 22894 6452
rect 14458 6372 14464 6384
rect 14108 6344 14464 6372
rect 14108 6316 14136 6344
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 17782 6375 17840 6381
rect 17782 6372 17794 6375
rect 16080 6344 17794 6372
rect 16080 6332 16086 6344
rect 17782 6341 17794 6344
rect 17828 6341 17840 6375
rect 18874 6372 18880 6384
rect 17782 6335 17840 6341
rect 18156 6344 18880 6372
rect 18156 6316 18184 6344
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 20162 6332 20168 6384
rect 20220 6372 20226 6384
rect 23106 6372 23112 6384
rect 20220 6344 23112 6372
rect 20220 6332 20226 6344
rect 13541 6307 13599 6313
rect 9548 6276 9996 6304
rect 9548 6264 9554 6276
rect 8386 6236 8392 6248
rect 8312 6208 8392 6236
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 9968 6236 9996 6276
rect 13541 6273 13553 6307
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 13814 6264 13820 6316
rect 13872 6264 13878 6316
rect 14090 6264 14096 6316
rect 14148 6264 14154 6316
rect 14349 6307 14407 6313
rect 14349 6304 14361 6307
rect 14200 6276 14361 6304
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 9968 6208 11529 6236
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 14200 6236 14228 6276
rect 14349 6273 14361 6276
rect 14395 6273 14407 6307
rect 14349 6267 14407 6273
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 18138 6304 18144 6316
rect 14700 6276 18144 6304
rect 14700 6264 14706 6276
rect 11517 6199 11575 6205
rect 13740 6208 14228 6236
rect 13740 6177 13768 6208
rect 15194 6196 15200 6248
rect 15252 6236 15258 6248
rect 16132 6245 16160 6276
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18506 6313 18512 6316
rect 18500 6267 18512 6313
rect 18506 6264 18512 6267
rect 18564 6264 18570 6316
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19961 6307 20019 6313
rect 19961 6304 19973 6307
rect 19024 6276 19973 6304
rect 19024 6264 19030 6276
rect 19961 6273 19973 6276
rect 20007 6273 20019 6307
rect 19961 6267 20019 6273
rect 21174 6264 21180 6316
rect 21232 6264 21238 6316
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6304 21511 6307
rect 21634 6304 21640 6316
rect 21499 6276 21640 6304
rect 21499 6273 21511 6276
rect 21453 6267 21511 6273
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 22756 6313 22784 6344
rect 23106 6332 23112 6344
rect 23164 6332 23170 6384
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6273 22799 6307
rect 22741 6267 22799 6273
rect 23658 6264 23664 6316
rect 23716 6264 23722 6316
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15252 6208 16037 6236
rect 15252 6196 15258 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6236 18107 6239
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 18095 6208 18245 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 19702 6236 19708 6248
rect 18233 6199 18291 6205
rect 19536 6208 19708 6236
rect 13725 6171 13783 6177
rect 13725 6137 13737 6171
rect 13771 6137 13783 6171
rect 13725 6131 13783 6137
rect 15470 6128 15476 6180
rect 15528 6128 15534 6180
rect 16040 6168 16068 6199
rect 16850 6168 16856 6180
rect 16040 6140 16856 6168
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 11287 6103 11345 6109
rect 11287 6100 11299 6103
rect 9732 6072 11299 6100
rect 9732 6060 9738 6072
rect 11287 6069 11299 6072
rect 11333 6069 11345 6103
rect 11287 6063 11345 6069
rect 13262 6060 13268 6112
rect 13320 6060 13326 6112
rect 13998 6060 14004 6112
rect 14056 6060 14062 6112
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 16942 6100 16948 6112
rect 16080 6072 16948 6100
rect 16080 6060 16086 6072
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18064 6100 18092 6199
rect 19536 6100 19564 6208
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 21542 6196 21548 6248
rect 21600 6236 21606 6248
rect 21600 6208 23520 6236
rect 21600 6196 21606 6208
rect 21085 6171 21143 6177
rect 21085 6137 21097 6171
rect 21131 6168 21143 6171
rect 21726 6168 21732 6180
rect 21131 6140 21732 6168
rect 21131 6137 21143 6140
rect 21085 6131 21143 6137
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 23492 6177 23520 6208
rect 23477 6171 23535 6177
rect 23477 6137 23489 6171
rect 23523 6137 23535 6171
rect 23477 6131 23535 6137
rect 17828 6072 19564 6100
rect 17828 6060 17834 6072
rect 22186 6060 22192 6112
rect 22244 6060 22250 6112
rect 1104 6010 24012 6032
rect 1104 5958 1350 6010
rect 1402 5958 1414 6010
rect 1466 5958 1478 6010
rect 1530 5958 1542 6010
rect 1594 5958 1606 6010
rect 1658 5958 4350 6010
rect 4402 5958 4414 6010
rect 4466 5958 4478 6010
rect 4530 5958 4542 6010
rect 4594 5958 4606 6010
rect 4658 5958 7350 6010
rect 7402 5958 7414 6010
rect 7466 5958 7478 6010
rect 7530 5958 7542 6010
rect 7594 5958 7606 6010
rect 7658 5958 10350 6010
rect 10402 5958 10414 6010
rect 10466 5958 10478 6010
rect 10530 5958 10542 6010
rect 10594 5958 10606 6010
rect 10658 5958 13350 6010
rect 13402 5958 13414 6010
rect 13466 5958 13478 6010
rect 13530 5958 13542 6010
rect 13594 5958 13606 6010
rect 13658 5958 16350 6010
rect 16402 5958 16414 6010
rect 16466 5958 16478 6010
rect 16530 5958 16542 6010
rect 16594 5958 16606 6010
rect 16658 5958 19350 6010
rect 19402 5958 19414 6010
rect 19466 5958 19478 6010
rect 19530 5958 19542 6010
rect 19594 5958 19606 6010
rect 19658 5958 22350 6010
rect 22402 5958 22414 6010
rect 22466 5958 22478 6010
rect 22530 5958 22542 6010
rect 22594 5958 22606 6010
rect 22658 5958 24012 6010
rect 1104 5936 24012 5958
rect 9766 5856 9772 5908
rect 9824 5856 9830 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 9916 5868 9965 5896
rect 9916 5856 9922 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 9953 5859 10011 5865
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12342 5896 12348 5908
rect 12299 5868 12348 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 15470 5856 15476 5908
rect 15528 5896 15534 5908
rect 15528 5868 16804 5896
rect 15528 5856 15534 5868
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5626 5760 5632 5772
rect 5123 5732 5632 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 12434 5760 12440 5772
rect 12406 5720 12440 5760
rect 12492 5720 12498 5772
rect 14090 5720 14096 5772
rect 14148 5720 14154 5772
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 16439 5763 16497 5769
rect 16439 5760 16451 5763
rect 15528 5732 16451 5760
rect 15528 5720 15534 5732
rect 16439 5729 16451 5732
rect 16485 5729 16497 5763
rect 16439 5723 16497 5729
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 16776 5760 16804 5868
rect 18506 5856 18512 5908
rect 18564 5856 18570 5908
rect 18966 5856 18972 5908
rect 19024 5856 19030 5908
rect 19886 5856 19892 5908
rect 19944 5856 19950 5908
rect 20809 5899 20867 5905
rect 20809 5865 20821 5899
rect 20855 5896 20867 5899
rect 21266 5896 21272 5908
rect 20855 5868 21272 5896
rect 20855 5865 20867 5868
rect 20809 5859 20867 5865
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 16853 5831 16911 5837
rect 16853 5797 16865 5831
rect 16899 5828 16911 5831
rect 16942 5828 16948 5840
rect 16899 5800 16948 5828
rect 16899 5797 16911 5800
rect 16853 5791 16911 5797
rect 16942 5788 16948 5800
rect 17000 5828 17006 5840
rect 19904 5828 19932 5856
rect 20438 5828 20444 5840
rect 17000 5800 20444 5828
rect 17000 5788 17006 5800
rect 20438 5788 20444 5800
rect 20496 5788 20502 5840
rect 22186 5828 22192 5840
rect 21284 5800 22192 5828
rect 16623 5732 16804 5760
rect 17313 5763 17371 5769
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 17313 5729 17325 5763
rect 17359 5760 17371 5763
rect 18230 5760 18236 5772
rect 17359 5732 18236 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 19702 5720 19708 5772
rect 19760 5760 19766 5772
rect 21284 5769 21312 5800
rect 22186 5788 22192 5800
rect 22244 5788 22250 5840
rect 19889 5763 19947 5769
rect 19889 5760 19901 5763
rect 19760 5732 19901 5760
rect 19760 5720 19766 5732
rect 19889 5729 19901 5732
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 21269 5763 21327 5769
rect 21269 5729 21281 5763
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 21499 5732 21680 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 6104 5664 6960 5692
rect 6104 5610 6132 5664
rect 6503 5627 6561 5633
rect 6503 5593 6515 5627
rect 6549 5624 6561 5627
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 6549 5596 6653 5624
rect 6549 5593 6561 5596
rect 6503 5587 6561 5593
rect 6641 5593 6653 5596
rect 6687 5624 6699 5627
rect 6730 5624 6736 5636
rect 6687 5596 6736 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 6822 5584 6828 5636
rect 6880 5584 6886 5636
rect 6932 5624 6960 5664
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 9122 5692 9128 5704
rect 7432 5664 9128 5692
rect 7432 5652 7438 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 9674 5692 9680 5704
rect 9539 5664 9680 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 7190 5624 7196 5636
rect 6932 5596 7196 5624
rect 7190 5584 7196 5596
rect 7248 5624 7254 5636
rect 8018 5624 8024 5636
rect 7248 5596 8024 5624
rect 7248 5584 7254 5596
rect 8018 5584 8024 5596
rect 8076 5584 8082 5636
rect 9416 5568 9444 5655
rect 9674 5652 9680 5664
rect 9732 5692 9738 5704
rect 9950 5692 9956 5704
rect 9732 5664 9956 5692
rect 9732 5652 9738 5664
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 10100 5664 10149 5692
rect 10100 5652 10106 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5692 12127 5695
rect 12406 5692 12434 5720
rect 12830 5695 12888 5701
rect 12830 5692 12842 5695
rect 12115 5664 12842 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 12830 5661 12842 5664
rect 12876 5661 12888 5695
rect 12830 5655 12888 5661
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14349 5695 14407 5701
rect 14349 5692 14361 5695
rect 14056 5664 14361 5692
rect 14056 5652 14062 5664
rect 14349 5661 14361 5664
rect 14395 5661 14407 5695
rect 14349 5655 14407 5661
rect 16298 5652 16304 5704
rect 16356 5652 16362 5704
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5692 17555 5695
rect 17586 5692 17592 5704
rect 17543 5664 17592 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18693 5695 18751 5701
rect 18693 5692 18705 5695
rect 18380 5664 18705 5692
rect 18380 5652 18386 5664
rect 18693 5661 18705 5664
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 21177 5695 21235 5701
rect 21177 5661 21189 5695
rect 21223 5692 21235 5695
rect 21542 5692 21548 5704
rect 21223 5664 21548 5692
rect 21223 5661 21235 5664
rect 21177 5655 21235 5661
rect 21542 5652 21548 5664
rect 21600 5652 21606 5704
rect 11514 5584 11520 5636
rect 11572 5584 11578 5636
rect 12437 5627 12495 5633
rect 12437 5593 12449 5627
rect 12483 5624 12495 5627
rect 12526 5624 12532 5636
rect 12483 5596 12532 5624
rect 12483 5593 12495 5596
rect 12437 5587 12495 5593
rect 7006 5516 7012 5568
rect 7064 5516 7070 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 12452 5556 12480 5587
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 12621 5627 12679 5633
rect 12621 5593 12633 5627
rect 12667 5624 12679 5627
rect 13262 5624 13268 5636
rect 12667 5596 13268 5624
rect 12667 5593 12679 5596
rect 12621 5587 12679 5593
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 20622 5584 20628 5636
rect 20680 5624 20686 5636
rect 21652 5624 21680 5732
rect 20680 5596 21680 5624
rect 20680 5584 20686 5596
rect 12759 5559 12817 5565
rect 12759 5556 12771 5559
rect 9456 5528 12771 5556
rect 9456 5516 9462 5528
rect 12759 5525 12771 5528
rect 12805 5525 12817 5559
rect 12759 5519 12817 5525
rect 15470 5516 15476 5568
rect 15528 5516 15534 5568
rect 15657 5559 15715 5565
rect 15657 5525 15669 5559
rect 15703 5556 15715 5559
rect 17678 5556 17684 5568
rect 15703 5528 17684 5556
rect 15703 5525 15715 5528
rect 15657 5519 15715 5525
rect 17678 5516 17684 5528
rect 17736 5516 17742 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21450 5556 21456 5568
rect 20772 5528 21456 5556
rect 20772 5516 20778 5528
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 1104 5466 24164 5488
rect 1104 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 3042 5466
rect 3094 5414 3106 5466
rect 3158 5414 5850 5466
rect 5902 5414 5914 5466
rect 5966 5414 5978 5466
rect 6030 5414 6042 5466
rect 6094 5414 6106 5466
rect 6158 5414 8850 5466
rect 8902 5414 8914 5466
rect 8966 5414 8978 5466
rect 9030 5414 9042 5466
rect 9094 5414 9106 5466
rect 9158 5414 11850 5466
rect 11902 5414 11914 5466
rect 11966 5414 11978 5466
rect 12030 5414 12042 5466
rect 12094 5414 12106 5466
rect 12158 5414 14850 5466
rect 14902 5414 14914 5466
rect 14966 5414 14978 5466
rect 15030 5414 15042 5466
rect 15094 5414 15106 5466
rect 15158 5414 17850 5466
rect 17902 5414 17914 5466
rect 17966 5414 17978 5466
rect 18030 5414 18042 5466
rect 18094 5414 18106 5466
rect 18158 5414 20850 5466
rect 20902 5414 20914 5466
rect 20966 5414 20978 5466
rect 21030 5414 21042 5466
rect 21094 5414 21106 5466
rect 21158 5414 23850 5466
rect 23902 5414 23914 5466
rect 23966 5414 23978 5466
rect 24030 5414 24042 5466
rect 24094 5414 24106 5466
rect 24158 5414 24164 5466
rect 1104 5392 24164 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 8662 5352 8668 5364
rect 6880 5324 8668 5352
rect 6880 5312 6886 5324
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 8938 5352 8944 5364
rect 8812 5324 8944 5352
rect 8812 5312 8818 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 15286 5312 15292 5364
rect 15344 5312 15350 5364
rect 16206 5312 16212 5364
rect 16264 5312 16270 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 16758 5352 16764 5364
rect 16715 5324 16764 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17494 5352 17500 5364
rect 17175 5324 17500 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 6730 5284 6736 5296
rect 5736 5256 6736 5284
rect 5736 5225 5764 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 5810 5108 5816 5160
rect 5868 5108 5874 5160
rect 6104 5148 6132 5179
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6840 5216 6868 5312
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 6696 5188 6868 5216
rect 6932 5256 7297 5284
rect 6696 5176 6702 5188
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 6104 5120 6377 5148
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5117 6791 5151
rect 6733 5111 6791 5117
rect 5629 5083 5687 5089
rect 5629 5049 5641 5083
rect 5675 5080 5687 5083
rect 6564 5080 6592 5111
rect 5675 5052 6592 5080
rect 6748 5080 6776 5111
rect 6822 5108 6828 5160
rect 6880 5108 6886 5160
rect 6932 5080 6960 5256
rect 7285 5253 7297 5256
rect 7331 5284 7343 5287
rect 7374 5284 7380 5296
rect 7331 5256 7380 5284
rect 7331 5253 7343 5256
rect 7285 5247 7343 5253
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 7926 5284 7932 5296
rect 7484 5256 7932 5284
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7484 5225 7512 5256
rect 7926 5244 7932 5256
rect 7984 5244 7990 5296
rect 8386 5284 8392 5296
rect 8036 5256 8392 5284
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5185 7159 5219
rect 7101 5179 7159 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 7742 5216 7748 5228
rect 7699 5188 7748 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7116 5148 7144 5179
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 8036 5225 8064 5256
rect 8386 5244 8392 5256
rect 8444 5284 8450 5296
rect 8846 5284 8852 5296
rect 8444 5256 8852 5284
rect 8444 5244 8450 5256
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 19978 5284 19984 5296
rect 19904 5256 19984 5284
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8570 5216 8576 5228
rect 8159 5188 8576 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8720 5188 8953 5216
rect 8720 5176 8726 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15528 5188 15853 5216
rect 15528 5176 15534 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 16393 5219 16451 5225
rect 16393 5216 16405 5219
rect 16172 5188 16405 5216
rect 16172 5176 16178 5188
rect 16393 5185 16405 5188
rect 16439 5185 16451 5219
rect 16393 5179 16451 5185
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16816 5188 17049 5216
rect 16816 5176 16822 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 19904 5216 19932 5256
rect 19978 5244 19984 5256
rect 20036 5244 20042 5296
rect 17037 5179 17095 5185
rect 17328 5188 19932 5216
rect 17328 5160 17356 5188
rect 7834 5148 7840 5160
rect 7116 5120 7840 5148
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 6748 5052 6960 5080
rect 5675 5049 5687 5052
rect 5629 5043 5687 5049
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7469 5083 7527 5089
rect 7469 5080 7481 5083
rect 7248 5052 7481 5080
rect 7248 5040 7254 5052
rect 7469 5049 7481 5052
rect 7515 5049 7527 5083
rect 7944 5080 7972 5111
rect 8202 5108 8208 5160
rect 8260 5108 8266 5160
rect 9214 5108 9220 5160
rect 9272 5108 9278 5160
rect 17310 5108 17316 5160
rect 17368 5108 17374 5160
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5148 18199 5151
rect 18230 5148 18236 5160
rect 18187 5120 18236 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 19904 5157 19932 5188
rect 20070 5176 20076 5228
rect 20128 5176 20134 5228
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 20027 5120 20545 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 8478 5080 8484 5092
rect 7944 5052 8484 5080
rect 7469 5043 7527 5049
rect 8478 5040 8484 5052
rect 8536 5080 8542 5092
rect 9398 5080 9404 5092
rect 8536 5052 9404 5080
rect 8536 5040 8542 5052
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 19702 5040 19708 5092
rect 19760 5080 19766 5092
rect 21100 5080 21128 5111
rect 19760 5052 21128 5080
rect 19760 5040 19766 5052
rect 5997 5015 6055 5021
rect 5997 4981 6009 5015
rect 6043 5012 6055 5015
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 6043 4984 7297 5012
rect 6043 4981 6055 4984
rect 5997 4975 6055 4981
rect 7285 4981 7297 4984
rect 7331 4981 7343 5015
rect 7285 4975 7343 4981
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 12342 5012 12348 5024
rect 8076 4984 12348 5012
rect 8076 4972 8082 4984
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 17494 4972 17500 5024
rect 17552 4972 17558 5024
rect 20441 5015 20499 5021
rect 20441 4981 20453 5015
rect 20487 5012 20499 5015
rect 21726 5012 21732 5024
rect 20487 4984 21732 5012
rect 20487 4981 20499 4984
rect 20441 4975 20499 4981
rect 21726 4972 21732 4984
rect 21784 4972 21790 5024
rect 1104 4922 24012 4944
rect 1104 4870 1350 4922
rect 1402 4870 1414 4922
rect 1466 4870 1478 4922
rect 1530 4870 1542 4922
rect 1594 4870 1606 4922
rect 1658 4870 4350 4922
rect 4402 4870 4414 4922
rect 4466 4870 4478 4922
rect 4530 4870 4542 4922
rect 4594 4870 4606 4922
rect 4658 4870 7350 4922
rect 7402 4870 7414 4922
rect 7466 4870 7478 4922
rect 7530 4870 7542 4922
rect 7594 4870 7606 4922
rect 7658 4870 10350 4922
rect 10402 4870 10414 4922
rect 10466 4870 10478 4922
rect 10530 4870 10542 4922
rect 10594 4870 10606 4922
rect 10658 4870 13350 4922
rect 13402 4870 13414 4922
rect 13466 4870 13478 4922
rect 13530 4870 13542 4922
rect 13594 4870 13606 4922
rect 13658 4870 16350 4922
rect 16402 4870 16414 4922
rect 16466 4870 16478 4922
rect 16530 4870 16542 4922
rect 16594 4870 16606 4922
rect 16658 4870 19350 4922
rect 19402 4870 19414 4922
rect 19466 4870 19478 4922
rect 19530 4870 19542 4922
rect 19594 4870 19606 4922
rect 19658 4870 22350 4922
rect 22402 4870 22414 4922
rect 22466 4870 22478 4922
rect 22530 4870 22542 4922
rect 22594 4870 22606 4922
rect 22658 4870 24012 4922
rect 1104 4848 24012 4870
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 8260 4780 9689 4808
rect 8260 4768 8266 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 9677 4771 9735 4777
rect 9861 4811 9919 4817
rect 9861 4777 9873 4811
rect 9907 4808 9919 4811
rect 11514 4808 11520 4820
rect 9907 4780 11520 4808
rect 9907 4777 9919 4780
rect 9861 4771 9919 4777
rect 7742 4740 7748 4752
rect 7116 4712 7748 4740
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 5868 4644 6561 4672
rect 5868 4632 5874 4644
rect 6549 4641 6561 4644
rect 6595 4672 6607 4675
rect 6914 4672 6920 4684
rect 6595 4644 6920 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7116 4681 7144 4712
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 9214 4700 9220 4752
rect 9272 4740 9278 4752
rect 9582 4740 9588 4752
rect 9272 4712 9588 4740
rect 9272 4700 9278 4712
rect 9582 4700 9588 4712
rect 9640 4740 9646 4752
rect 9876 4740 9904 4771
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 9640 4712 9904 4740
rect 9640 4700 9646 4712
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7190 4632 7196 4684
rect 7248 4632 7254 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7892 4644 8033 4672
rect 7892 4632 7898 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8662 4672 8668 4684
rect 8021 4635 8079 4641
rect 8220 4644 8668 4672
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 6822 4604 6828 4616
rect 6411 4576 6828 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 8220 4613 8248 4644
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 8846 4632 8852 4684
rect 8904 4632 8910 4684
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9232 4672 9260 4700
rect 9426 4675 9484 4681
rect 9426 4672 9438 4675
rect 8987 4644 9260 4672
rect 9324 4644 9438 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 8864 4604 8892 4632
rect 9324 4604 9352 4644
rect 9426 4641 9438 4644
rect 9472 4672 9484 4675
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 9472 4644 10241 4672
rect 9472 4641 9484 4644
rect 9426 4635 9484 4641
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10229 4635 10287 4641
rect 15654 4632 15660 4684
rect 15712 4632 15718 4684
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 18417 4675 18475 4681
rect 18417 4672 18429 4675
rect 18380 4644 18429 4672
rect 18380 4632 18386 4644
rect 18417 4641 18429 4644
rect 18463 4641 18475 4675
rect 18417 4635 18475 4641
rect 18601 4675 18659 4681
rect 18601 4641 18613 4675
rect 18647 4672 18659 4675
rect 19794 4672 19800 4684
rect 18647 4644 19800 4672
rect 18647 4641 18659 4644
rect 18601 4635 18659 4641
rect 19794 4632 19800 4644
rect 19852 4672 19858 4684
rect 20070 4672 20076 4684
rect 19852 4644 20076 4672
rect 19852 4632 19858 4644
rect 20070 4632 20076 4644
rect 20128 4632 20134 4684
rect 8864 4576 9352 4604
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10781 4607 10839 4613
rect 9640 4576 9904 4604
rect 9640 4564 9646 4576
rect 7837 4539 7895 4545
rect 7837 4505 7849 4539
rect 7883 4536 7895 4539
rect 7926 4536 7932 4548
rect 7883 4508 7932 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 9876 4545 9904 4576
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 8628 4508 9321 4536
rect 8628 4496 8634 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9309 4499 9367 4505
rect 9861 4539 9919 4545
rect 9861 4505 9873 4539
rect 9907 4505 9919 4539
rect 10796 4536 10824 4567
rect 10870 4564 10876 4616
rect 10928 4564 10934 4616
rect 12342 4564 12348 4616
rect 12400 4564 12406 4616
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 19978 4604 19984 4616
rect 19935 4576 19984 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 10962 4536 10968 4548
rect 10796 4508 10968 4536
rect 9861 4499 9919 4505
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 15924 4539 15982 4545
rect 15924 4505 15936 4539
rect 15970 4536 15982 4539
rect 16850 4536 16856 4548
rect 15970 4508 16856 4536
rect 15970 4505 15982 4508
rect 15924 4499 15982 4505
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 17129 4539 17187 4545
rect 17129 4536 17141 4539
rect 17000 4508 17141 4536
rect 17000 4496 17006 4508
rect 17129 4505 17141 4508
rect 17175 4505 17187 4539
rect 17129 4499 17187 4505
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5776 4440 5917 4468
rect 5776 4428 5782 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 5905 4431 5963 4437
rect 6270 4428 6276 4480
rect 6328 4428 6334 4480
rect 7282 4428 7288 4480
rect 7340 4428 7346 4480
rect 7653 4471 7711 4477
rect 7653 4437 7665 4471
rect 7699 4468 7711 4471
rect 7742 4468 7748 4480
rect 7699 4440 7748 4468
rect 7699 4437 7711 4440
rect 7653 4431 7711 4437
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 7944 4468 7972 4496
rect 9214 4468 9220 4480
rect 7944 4440 9220 4468
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9582 4428 9588 4480
rect 9640 4428 9646 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 10778 4468 10784 4480
rect 10643 4440 10784 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 12308 4440 12449 4468
rect 12308 4428 12314 4440
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 17034 4428 17040 4480
rect 17092 4468 17098 4480
rect 17696 4468 17724 4567
rect 19978 4564 19984 4576
rect 20036 4604 20042 4616
rect 20254 4604 20260 4616
rect 20036 4576 20260 4604
rect 20036 4564 20042 4576
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 21358 4564 21364 4616
rect 21416 4564 21422 4616
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 19245 4539 19303 4545
rect 19245 4536 19257 4539
rect 18739 4508 19257 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 19245 4505 19257 4508
rect 19291 4505 19303 4539
rect 19245 4499 19303 4505
rect 21116 4539 21174 4545
rect 21116 4505 21128 4539
rect 21162 4536 21174 4539
rect 21266 4536 21272 4548
rect 21162 4508 21272 4536
rect 21162 4505 21174 4508
rect 21116 4499 21174 4505
rect 21266 4496 21272 4508
rect 21324 4496 21330 4548
rect 17092 4440 17724 4468
rect 17092 4428 17098 4440
rect 18874 4428 18880 4480
rect 18932 4468 18938 4480
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 18932 4440 19073 4468
rect 18932 4428 18938 4440
rect 19061 4437 19073 4440
rect 19107 4437 19119 4471
rect 19061 4431 19119 4437
rect 19518 4428 19524 4480
rect 19576 4468 19582 4480
rect 19981 4471 20039 4477
rect 19981 4468 19993 4471
rect 19576 4440 19993 4468
rect 19576 4428 19582 4440
rect 19981 4437 19993 4440
rect 20027 4468 20039 4471
rect 20070 4468 20076 4480
rect 20027 4440 20076 4468
rect 20027 4437 20039 4440
rect 19981 4431 20039 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 1104 4378 24164 4400
rect 1104 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 3042 4378
rect 3094 4326 3106 4378
rect 3158 4326 5850 4378
rect 5902 4326 5914 4378
rect 5966 4326 5978 4378
rect 6030 4326 6042 4378
rect 6094 4326 6106 4378
rect 6158 4326 8850 4378
rect 8902 4326 8914 4378
rect 8966 4326 8978 4378
rect 9030 4326 9042 4378
rect 9094 4326 9106 4378
rect 9158 4326 11850 4378
rect 11902 4326 11914 4378
rect 11966 4326 11978 4378
rect 12030 4326 12042 4378
rect 12094 4326 12106 4378
rect 12158 4326 14850 4378
rect 14902 4326 14914 4378
rect 14966 4326 14978 4378
rect 15030 4326 15042 4378
rect 15094 4326 15106 4378
rect 15158 4326 17850 4378
rect 17902 4326 17914 4378
rect 17966 4326 17978 4378
rect 18030 4326 18042 4378
rect 18094 4326 18106 4378
rect 18158 4326 20850 4378
rect 20902 4326 20914 4378
rect 20966 4326 20978 4378
rect 21030 4326 21042 4378
rect 21094 4326 21106 4378
rect 21158 4326 23850 4378
rect 23902 4326 23914 4378
rect 23966 4326 23978 4378
rect 24030 4326 24042 4378
rect 24094 4326 24106 4378
rect 24158 4326 24164 4378
rect 1104 4304 24164 4326
rect 6457 4267 6515 4273
rect 6457 4233 6469 4267
rect 6503 4264 6515 4267
rect 6822 4264 6828 4276
rect 6503 4236 6828 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7469 4267 7527 4273
rect 7469 4264 7481 4267
rect 7340 4236 7481 4264
rect 7340 4224 7346 4236
rect 7469 4233 7481 4236
rect 7515 4233 7527 4267
rect 9398 4264 9404 4276
rect 7469 4227 7527 4233
rect 8496 4236 9404 4264
rect 8496 4140 8524 4236
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 10226 4224 10232 4276
rect 10284 4264 10290 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10284 4236 10517 4264
rect 10284 4224 10290 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10505 4227 10563 4233
rect 17129 4267 17187 4273
rect 17129 4233 17141 4267
rect 17175 4264 17187 4267
rect 17494 4264 17500 4276
rect 17175 4236 17500 4264
rect 17175 4233 17187 4236
rect 17129 4227 17187 4233
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 19153 4267 19211 4273
rect 19153 4233 19165 4267
rect 19199 4264 19211 4267
rect 20346 4264 20352 4276
rect 19199 4236 20352 4264
rect 19199 4233 19211 4236
rect 19153 4227 19211 4233
rect 20346 4224 20352 4236
rect 20404 4224 20410 4276
rect 21266 4224 21272 4276
rect 21324 4224 21330 4276
rect 8757 4199 8815 4205
rect 8757 4165 8769 4199
rect 8803 4196 8815 4199
rect 8803 4168 9812 4196
rect 8803 4165 8815 4168
rect 8757 4159 8815 4165
rect 5718 4088 5724 4140
rect 5776 4088 5782 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 6328 4100 6377 4128
rect 6328 4088 6334 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6638 4128 6644 4140
rect 6595 4100 6644 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6380 4060 6408 4091
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 7926 4128 7932 4140
rect 7699 4100 7932 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 7926 4088 7932 4100
rect 7984 4128 7990 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 7984 4100 8033 4128
rect 7984 4088 7990 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8478 4088 8484 4140
rect 8536 4088 8542 4140
rect 6822 4060 6828 4072
rect 6380 4032 6828 4060
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 6972 4032 7849 4060
rect 6972 4020 6978 4032
rect 7837 4029 7849 4032
rect 7883 4060 7895 4063
rect 8202 4060 8208 4072
rect 7883 4032 8208 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8772 4060 8800 4159
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9398 4128 9404 4140
rect 9263 4100 9404 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 9784 4128 9812 4168
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 11149 4199 11207 4205
rect 11149 4196 11161 4199
rect 10928 4168 11161 4196
rect 10928 4156 10934 4168
rect 11149 4165 11161 4168
rect 11195 4165 11207 4199
rect 11149 4159 11207 4165
rect 12250 4156 12256 4208
rect 12308 4156 12314 4208
rect 13814 4196 13820 4208
rect 13648 4168 13820 4196
rect 9784 4100 11008 4128
rect 10980 4072 11008 4100
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 11698 4128 11704 4140
rect 11388 4100 11704 4128
rect 11388 4088 11394 4100
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13311 4100 13461 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13449 4097 13461 4100
rect 13495 4128 13507 4131
rect 13648 4128 13676 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 16206 4156 16212 4208
rect 16264 4156 16270 4208
rect 13722 4137 13728 4140
rect 13495 4100 13676 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13716 4091 13728 4137
rect 13722 4088 13728 4091
rect 13780 4088 13786 4140
rect 13832 4128 13860 4156
rect 15654 4128 15660 4140
rect 13832 4100 15660 4128
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16224 4128 16252 4156
rect 17037 4131 17095 4137
rect 15988 4100 16804 4128
rect 15988 4088 15994 4100
rect 8496 4032 8800 4060
rect 9125 4063 9183 4069
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8496 3933 8524 4032
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9766 4060 9772 4072
rect 9171 4032 9772 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10686 4060 10692 4072
rect 10428 4032 10692 4060
rect 8665 3995 8723 4001
rect 8665 3961 8677 3995
rect 8711 3992 8723 3995
rect 8754 3992 8760 4004
rect 8711 3964 8760 3992
rect 8711 3961 8723 3964
rect 8665 3955 8723 3961
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 9306 3952 9312 4004
rect 9364 3992 9370 4004
rect 9401 3995 9459 4001
rect 9401 3992 9413 3995
rect 9364 3964 9413 3992
rect 9364 3952 9370 3964
rect 9401 3961 9413 3964
rect 9447 3961 9459 3995
rect 9401 3955 9459 3961
rect 9858 3952 9864 4004
rect 9916 3952 9922 4004
rect 10428 4001 10456 4032
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11020 4032 11529 4060
rect 11020 4020 11026 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 12986 4020 12992 4072
rect 13044 4020 13050 4072
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 14792 4032 15485 4060
rect 14792 4020 14798 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3961 10471 3995
rect 10413 3955 10471 3961
rect 10597 3995 10655 4001
rect 10597 3961 10609 3995
rect 10643 3992 10655 3995
rect 10870 3992 10876 4004
rect 10643 3964 10876 3992
rect 10643 3961 10655 3964
rect 10597 3955 10655 3961
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 14829 3995 14887 4001
rect 14829 3961 14841 3995
rect 14875 3992 14887 3995
rect 16114 3992 16120 4004
rect 14875 3964 16120 3992
rect 14875 3961 14887 3964
rect 14829 3955 14887 3961
rect 16114 3952 16120 3964
rect 16172 3992 16178 4004
rect 16224 3992 16252 4023
rect 16172 3964 16252 3992
rect 16172 3952 16178 3964
rect 8481 3927 8539 3933
rect 8481 3924 8493 3927
rect 8352 3896 8493 3924
rect 8352 3884 8358 3896
rect 8481 3893 8493 3896
rect 8527 3893 8539 3927
rect 8481 3887 8539 3893
rect 9214 3884 9220 3936
rect 9272 3884 9278 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9548 3896 10241 3924
rect 9548 3884 9554 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 14918 3884 14924 3936
rect 14976 3884 14982 3936
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15436 3896 15669 3924
rect 15436 3884 15442 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 15746 3884 15752 3936
rect 15804 3924 15810 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 15804 3896 16681 3924
rect 15804 3884 15810 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16776 3924 16804 4100
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17126 4128 17132 4140
rect 17083 4100 17132 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17460 4100 17693 4128
rect 17460 4088 17466 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 18040 4131 18098 4137
rect 18040 4097 18052 4131
rect 18086 4128 18098 4131
rect 18322 4128 18328 4140
rect 18086 4100 18328 4128
rect 18086 4097 18098 4100
rect 18040 4091 18098 4097
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 19337 4131 19395 4137
rect 19337 4097 19349 4131
rect 19383 4128 19395 4131
rect 19702 4128 19708 4140
rect 19383 4100 19708 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 20254 4088 20260 4140
rect 20312 4088 20318 4140
rect 20346 4088 20352 4140
rect 20404 4137 20410 4140
rect 20404 4131 20432 4137
rect 20420 4097 20432 4131
rect 20404 4091 20432 4097
rect 20404 4088 20410 4091
rect 21450 4088 21456 4140
rect 21508 4088 21514 4140
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 17770 4020 17776 4072
rect 17828 4020 17834 4072
rect 19518 4020 19524 4072
rect 19576 4020 19582 4072
rect 20533 4063 20591 4069
rect 20533 4060 20545 4063
rect 19628 4032 20545 4060
rect 16850 3952 16856 4004
rect 16908 3992 16914 4004
rect 17497 3995 17555 4001
rect 17497 3992 17509 3995
rect 16908 3964 17509 3992
rect 16908 3952 16914 3964
rect 17497 3961 17509 3964
rect 17543 3961 17555 3995
rect 17497 3955 17555 3961
rect 19628 3924 19656 4032
rect 20533 4029 20545 4032
rect 20579 4060 20591 4063
rect 20714 4060 20720 4072
rect 20579 4032 20720 4060
rect 20579 4029 20591 4032
rect 20533 4023 20591 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 22066 4032 22385 4060
rect 19886 3952 19892 4004
rect 19944 3992 19950 4004
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 19944 3964 19993 3992
rect 19944 3952 19950 3964
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 22066 3992 22094 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 19981 3955 20039 3961
rect 20916 3964 22094 3992
rect 16776 3896 19656 3924
rect 16669 3887 16727 3893
rect 20070 3884 20076 3936
rect 20128 3924 20134 3936
rect 20916 3924 20944 3964
rect 20128 3896 20944 3924
rect 21177 3927 21235 3933
rect 20128 3884 20134 3896
rect 21177 3893 21189 3927
rect 21223 3924 21235 3927
rect 21634 3924 21640 3936
rect 21223 3896 21640 3924
rect 21223 3893 21235 3896
rect 21177 3887 21235 3893
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 21818 3884 21824 3936
rect 21876 3884 21882 3936
rect 1104 3834 24012 3856
rect 1104 3782 1350 3834
rect 1402 3782 1414 3834
rect 1466 3782 1478 3834
rect 1530 3782 1542 3834
rect 1594 3782 1606 3834
rect 1658 3782 4350 3834
rect 4402 3782 4414 3834
rect 4466 3782 4478 3834
rect 4530 3782 4542 3834
rect 4594 3782 4606 3834
rect 4658 3782 7350 3834
rect 7402 3782 7414 3834
rect 7466 3782 7478 3834
rect 7530 3782 7542 3834
rect 7594 3782 7606 3834
rect 7658 3782 10350 3834
rect 10402 3782 10414 3834
rect 10466 3782 10478 3834
rect 10530 3782 10542 3834
rect 10594 3782 10606 3834
rect 10658 3782 13350 3834
rect 13402 3782 13414 3834
rect 13466 3782 13478 3834
rect 13530 3782 13542 3834
rect 13594 3782 13606 3834
rect 13658 3782 16350 3834
rect 16402 3782 16414 3834
rect 16466 3782 16478 3834
rect 16530 3782 16542 3834
rect 16594 3782 16606 3834
rect 16658 3782 19350 3834
rect 19402 3782 19414 3834
rect 19466 3782 19478 3834
rect 19530 3782 19542 3834
rect 19594 3782 19606 3834
rect 19658 3782 22350 3834
rect 22402 3782 22414 3834
rect 22466 3782 22478 3834
rect 22530 3782 22542 3834
rect 22594 3782 22606 3834
rect 22658 3782 24012 3834
rect 1104 3760 24012 3782
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 9030 3720 9036 3732
rect 8444 3692 9036 3720
rect 8444 3680 8450 3692
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9125 3723 9183 3729
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 9214 3720 9220 3732
rect 9171 3692 9220 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10226 3720 10232 3732
rect 9907 3692 10232 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10836 3692 11161 3720
rect 10836 3680 10842 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 13780 3692 15025 3720
rect 13780 3680 13786 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 17221 3723 17279 3729
rect 16080 3692 16528 3720
rect 16080 3680 16086 3692
rect 7377 3655 7435 3661
rect 7377 3652 7389 3655
rect 6656 3624 7389 3652
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 4764 3556 5273 3584
rect 4764 3544 4770 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 5534 3544 5540 3596
rect 5592 3544 5598 3596
rect 6656 3502 6684 3624
rect 7377 3621 7389 3624
rect 7423 3652 7435 3655
rect 7926 3652 7932 3664
rect 7423 3624 7932 3652
rect 7423 3621 7435 3624
rect 7377 3615 7435 3621
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8662 3652 8668 3664
rect 8076 3624 8668 3652
rect 8076 3612 8082 3624
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 9490 3652 9496 3664
rect 9232 3624 9496 3652
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6880 3556 7021 3584
rect 6880 3544 6886 3556
rect 7009 3553 7021 3556
rect 7055 3584 7067 3587
rect 8294 3584 8300 3596
rect 7055 3556 8300 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8536 3556 8585 3584
rect 8536 3544 8542 3556
rect 8573 3553 8585 3556
rect 8619 3553 8631 3587
rect 8573 3547 8631 3553
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 9232 3584 9260 3624
rect 9490 3612 9496 3624
rect 9548 3612 9554 3664
rect 9766 3612 9772 3664
rect 9824 3652 9830 3664
rect 16500 3661 16528 3692
rect 17221 3689 17233 3723
rect 17267 3720 17279 3723
rect 18230 3720 18236 3732
rect 17267 3692 18236 3720
rect 17267 3689 17279 3692
rect 17221 3683 17279 3689
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 9824 3624 11713 3652
rect 9824 3612 9830 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 11701 3615 11759 3621
rect 14185 3655 14243 3661
rect 14185 3621 14197 3655
rect 14231 3621 14243 3655
rect 14185 3615 14243 3621
rect 16485 3655 16543 3661
rect 16485 3621 16497 3655
rect 16531 3621 16543 3655
rect 16485 3615 16543 3621
rect 8803 3556 9260 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 7742 3516 7748 3528
rect 7699 3488 7748 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8386 3516 8392 3528
rect 8036 3488 8392 3516
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 7282 3448 7288 3460
rect 7239 3420 7288 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 8036 3457 8064 3488
rect 8386 3476 8392 3488
rect 8444 3516 8450 3528
rect 9232 3525 9260 3556
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3584 9367 3587
rect 10229 3587 10287 3593
rect 10229 3584 10241 3587
rect 9355 3556 10241 3584
rect 9355 3553 9367 3556
rect 9309 3547 9367 3553
rect 10229 3553 10241 3556
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 10778 3584 10784 3596
rect 10468 3556 10784 3584
rect 10468 3544 10474 3556
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 13449 3587 13507 3593
rect 13449 3553 13461 3587
rect 13495 3584 13507 3587
rect 13814 3584 13820 3596
rect 13495 3556 13820 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8444 3488 8953 3516
rect 8444 3476 8450 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9582 3516 9588 3528
rect 9447 3488 9588 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 9582 3476 9588 3488
rect 9640 3516 9646 3528
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 9640 3488 11529 3516
rect 9640 3476 9646 3488
rect 11517 3485 11529 3488
rect 11563 3485 11575 3519
rect 11517 3479 11575 3485
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 14200 3516 14228 3615
rect 14642 3544 14648 3596
rect 14700 3584 14706 3596
rect 16114 3593 16120 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14700 3556 14749 3584
rect 14700 3544 14706 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 16092 3587 16120 3593
rect 16092 3553 16104 3587
rect 16092 3547 16120 3553
rect 16114 3544 16120 3547
rect 16172 3544 16178 3596
rect 16945 3587 17003 3593
rect 16945 3553 16957 3587
rect 16991 3584 17003 3587
rect 17034 3584 17040 3596
rect 16991 3556 17040 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 17236 3584 17264 3683
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 19429 3723 19487 3729
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 19702 3720 19708 3732
rect 19475 3692 19708 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 20438 3680 20444 3732
rect 20496 3720 20502 3732
rect 20496 3692 21404 3720
rect 20496 3680 20502 3692
rect 21376 3652 21404 3692
rect 21376 3624 21496 3652
rect 17175 3556 17264 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 13955 3488 14228 3516
rect 14553 3519 14611 3525
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 14553 3485 14565 3519
rect 14599 3516 14611 3519
rect 14918 3516 14924 3528
rect 14599 3488 14924 3516
rect 14599 3485 14611 3488
rect 14553 3479 14611 3485
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 15194 3476 15200 3528
rect 15252 3476 15258 3528
rect 15286 3476 15292 3528
rect 15344 3476 15350 3528
rect 15930 3476 15936 3528
rect 15988 3476 15994 3528
rect 16206 3476 16212 3528
rect 16264 3476 16270 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 17828 3488 18613 3516
rect 17828 3476 17834 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 8021 3451 8079 3457
rect 8021 3417 8033 3451
rect 8067 3417 8079 3451
rect 8021 3411 8079 3417
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9490 3448 9496 3460
rect 9088 3420 9496 3448
rect 9088 3408 9094 3420
rect 9490 3408 9496 3420
rect 9548 3448 9554 3460
rect 9858 3448 9864 3460
rect 9548 3420 9864 3448
rect 9548 3408 9554 3420
rect 9858 3408 9864 3420
rect 9916 3448 9922 3460
rect 9916 3420 10180 3448
rect 9916 3408 9922 3420
rect 7469 3383 7527 3389
rect 7469 3349 7481 3383
rect 7515 3380 7527 3383
rect 7558 3380 7564 3392
rect 7515 3352 7564 3380
rect 7515 3349 7527 3352
rect 7469 3343 7527 3349
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8481 3383 8539 3389
rect 8481 3380 8493 3383
rect 8352 3352 8493 3380
rect 8352 3340 8358 3352
rect 8481 3349 8493 3352
rect 8527 3380 8539 3383
rect 9398 3380 9404 3392
rect 8527 3352 9404 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 10042 3340 10048 3392
rect 10100 3340 10106 3392
rect 10152 3380 10180 3420
rect 10226 3408 10232 3460
rect 10284 3448 10290 3460
rect 10505 3451 10563 3457
rect 10505 3448 10517 3451
rect 10284 3420 10517 3448
rect 10284 3408 10290 3420
rect 10505 3417 10517 3420
rect 10551 3417 10563 3451
rect 11149 3451 11207 3457
rect 11149 3448 11161 3451
rect 10505 3411 10563 3417
rect 10612 3420 11161 3448
rect 10612 3380 10640 3420
rect 11149 3417 11161 3420
rect 11195 3417 11207 3451
rect 11149 3411 11207 3417
rect 12158 3408 12164 3460
rect 12216 3408 12222 3460
rect 13170 3408 13176 3460
rect 13228 3408 13234 3460
rect 14645 3451 14703 3457
rect 14645 3417 14657 3451
rect 14691 3448 14703 3451
rect 15304 3448 15332 3476
rect 14691 3420 15332 3448
rect 14691 3417 14703 3420
rect 14645 3411 14703 3417
rect 17310 3408 17316 3460
rect 17368 3448 17374 3460
rect 18334 3451 18392 3457
rect 18334 3448 18346 3451
rect 17368 3420 18346 3448
rect 17368 3408 17374 3420
rect 18334 3417 18346 3420
rect 18380 3417 18392 3451
rect 18616 3448 18644 3479
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 19628 3488 20821 3516
rect 19628 3448 19656 3488
rect 20809 3485 20821 3488
rect 20855 3516 20867 3519
rect 21358 3516 21364 3528
rect 20855 3488 21364 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21468 3525 21496 3624
rect 21634 3544 21640 3596
rect 21692 3584 21698 3596
rect 21692 3556 22140 3584
rect 21692 3544 21698 3556
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 21726 3476 21732 3528
rect 21784 3516 21790 3528
rect 22112 3525 22140 3556
rect 21821 3519 21879 3525
rect 21821 3516 21833 3519
rect 21784 3488 21833 3516
rect 21784 3476 21790 3488
rect 21821 3485 21833 3488
rect 21867 3485 21879 3519
rect 21821 3479 21879 3485
rect 22097 3519 22155 3525
rect 22097 3485 22109 3519
rect 22143 3485 22155 3519
rect 22097 3479 22155 3485
rect 18616 3420 19656 3448
rect 20564 3451 20622 3457
rect 18334 3411 18392 3417
rect 20564 3417 20576 3451
rect 20610 3448 20622 3451
rect 20610 3420 21680 3448
rect 20610 3417 20622 3420
rect 20564 3411 20622 3417
rect 10152 3352 10640 3380
rect 10870 3340 10876 3392
rect 10928 3340 10934 3392
rect 10962 3340 10968 3392
rect 11020 3340 11026 3392
rect 13722 3340 13728 3392
rect 13780 3340 13786 3392
rect 15289 3383 15347 3389
rect 15289 3349 15301 3383
rect 15335 3380 15347 3383
rect 17126 3380 17132 3392
rect 15335 3352 17132 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 18690 3340 18696 3392
rect 18748 3340 18754 3392
rect 19702 3340 19708 3392
rect 19760 3380 19766 3392
rect 21652 3389 21680 3420
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 19760 3352 20913 3380
rect 19760 3340 19766 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 21637 3383 21695 3389
rect 21637 3349 21649 3383
rect 21683 3349 21695 3383
rect 21637 3343 21695 3349
rect 21910 3340 21916 3392
rect 21968 3340 21974 3392
rect 1104 3290 24164 3312
rect 1104 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 3042 3290
rect 3094 3238 3106 3290
rect 3158 3238 5850 3290
rect 5902 3238 5914 3290
rect 5966 3238 5978 3290
rect 6030 3238 6042 3290
rect 6094 3238 6106 3290
rect 6158 3238 8850 3290
rect 8902 3238 8914 3290
rect 8966 3238 8978 3290
rect 9030 3238 9042 3290
rect 9094 3238 9106 3290
rect 9158 3238 11850 3290
rect 11902 3238 11914 3290
rect 11966 3238 11978 3290
rect 12030 3238 12042 3290
rect 12094 3238 12106 3290
rect 12158 3238 14850 3290
rect 14902 3238 14914 3290
rect 14966 3238 14978 3290
rect 15030 3238 15042 3290
rect 15094 3238 15106 3290
rect 15158 3238 17850 3290
rect 17902 3238 17914 3290
rect 17966 3238 17978 3290
rect 18030 3238 18042 3290
rect 18094 3238 18106 3290
rect 18158 3238 20850 3290
rect 20902 3238 20914 3290
rect 20966 3238 20978 3290
rect 21030 3238 21042 3290
rect 21094 3238 21106 3290
rect 21158 3238 23850 3290
rect 23902 3238 23914 3290
rect 23966 3238 23978 3290
rect 24030 3238 24042 3290
rect 24094 3238 24106 3290
rect 24158 3238 24164 3290
rect 1104 3216 24164 3238
rect 7558 3176 7564 3188
rect 6932 3148 7564 3176
rect 6932 3117 6960 3148
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 8386 3136 8392 3188
rect 8444 3136 8450 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 9548 3148 9597 3176
rect 9548 3136 9554 3148
rect 9585 3145 9597 3148
rect 9631 3145 9643 3179
rect 9585 3139 9643 3145
rect 10410 3136 10416 3188
rect 10468 3136 10474 3188
rect 11330 3176 11336 3188
rect 10520 3148 11336 3176
rect 6917 3111 6975 3117
rect 6917 3077 6929 3111
rect 6963 3077 6975 3111
rect 6917 3071 6975 3077
rect 7926 3068 7932 3120
rect 7984 3068 7990 3120
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 10520 3108 10548 3148
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11701 3179 11759 3185
rect 11701 3145 11713 3179
rect 11747 3176 11759 3179
rect 13170 3176 13176 3188
rect 11747 3148 13176 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 14829 3179 14887 3185
rect 14829 3176 14841 3179
rect 14792 3148 14841 3176
rect 14792 3136 14798 3148
rect 14829 3145 14841 3148
rect 14875 3145 14887 3179
rect 14829 3139 14887 3145
rect 14921 3179 14979 3185
rect 14921 3145 14933 3179
rect 14967 3176 14979 3179
rect 15194 3176 15200 3188
rect 14967 3148 15200 3176
rect 14967 3145 14979 3148
rect 14921 3139 14979 3145
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 15378 3136 15384 3188
rect 15436 3136 15442 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3145 15991 3179
rect 15933 3139 15991 3145
rect 8260 3080 10548 3108
rect 8260 3068 8266 3080
rect 10686 3068 10692 3120
rect 10744 3068 10750 3120
rect 13814 3108 13820 3120
rect 13464 3080 13820 3108
rect 6178 3000 6184 3052
rect 6236 3040 6242 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 6236 3012 6653 3040
rect 6236 3000 6242 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10100 3012 10885 3040
rect 10100 3000 10106 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10962 3000 10968 3052
rect 11020 3000 11026 3052
rect 13464 3049 13492 3080
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15948 3108 15976 3139
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17034 3136 17040 3188
rect 17092 3136 17098 3188
rect 17402 3136 17408 3188
rect 17460 3136 17466 3188
rect 19702 3136 19708 3188
rect 19760 3136 19766 3188
rect 20441 3179 20499 3185
rect 20441 3176 20453 3179
rect 19812 3148 20453 3176
rect 19812 3120 19840 3148
rect 20441 3145 20453 3148
rect 20487 3145 20499 3179
rect 20441 3139 20499 3145
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3176 20867 3179
rect 21450 3176 21456 3188
rect 20855 3148 21456 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 21450 3136 21456 3148
rect 21508 3136 21514 3188
rect 17310 3108 17316 3120
rect 15344 3080 15884 3108
rect 15948 3080 17316 3108
rect 15344 3068 15350 3080
rect 13722 3049 13728 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11164 3012 11529 3040
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 10226 2972 10232 2984
rect 9640 2944 10232 2972
rect 9640 2932 9646 2944
rect 10226 2932 10232 2944
rect 10284 2932 10290 2984
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 11164 2913 11192 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13716 3040 13728 3049
rect 13683 3012 13728 3040
rect 13449 3003 13507 3009
rect 13716 3003 13728 3012
rect 13722 3000 13728 3003
rect 13780 3000 13786 3052
rect 15746 3000 15752 3052
rect 15804 3000 15810 3052
rect 15856 3040 15884 3080
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 18040 3111 18098 3117
rect 18040 3077 18052 3111
rect 18086 3108 18098 3111
rect 18690 3108 18696 3120
rect 18086 3080 18696 3108
rect 18086 3077 18098 3080
rect 18040 3071 18098 3077
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 19794 3108 19800 3120
rect 19659 3080 19800 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 20349 3111 20407 3117
rect 20349 3077 20361 3111
rect 20395 3108 20407 3111
rect 21818 3108 21824 3120
rect 20395 3080 21824 3108
rect 20395 3077 20407 3080
rect 20349 3071 20407 3077
rect 21818 3068 21824 3080
rect 21876 3068 21882 3120
rect 17034 3040 17040 3052
rect 15856 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 17184 3012 17693 3040
rect 17184 3000 17190 3012
rect 17681 3009 17693 3012
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 17770 3000 17776 3052
rect 17828 3000 17834 3052
rect 20622 3040 20628 3052
rect 17880 3012 20628 3040
rect 15562 2932 15568 2984
rect 15620 2932 15626 2984
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2972 16911 2975
rect 17218 2972 17224 2984
rect 16899 2944 17224 2972
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 17218 2932 17224 2944
rect 17276 2972 17282 2984
rect 17880 2972 17908 3012
rect 20180 2981 20208 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 17276 2944 17908 2972
rect 18800 2944 19809 2972
rect 17276 2932 17282 2944
rect 10045 2907 10103 2913
rect 10045 2904 10057 2907
rect 9548 2876 10057 2904
rect 9548 2864 9554 2876
rect 10045 2873 10057 2876
rect 10091 2873 10103 2907
rect 10045 2867 10103 2873
rect 11149 2907 11207 2913
rect 11149 2873 11161 2907
rect 11195 2873 11207 2907
rect 15580 2904 15608 2932
rect 15580 2876 17632 2904
rect 11149 2867 11207 2873
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 10134 2836 10140 2848
rect 7340 2808 10140 2836
rect 7340 2796 7346 2808
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 10597 2839 10655 2845
rect 10597 2805 10609 2839
rect 10643 2836 10655 2839
rect 10689 2839 10747 2845
rect 10689 2836 10701 2839
rect 10643 2808 10701 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 10689 2805 10701 2808
rect 10735 2805 10747 2839
rect 10689 2799 10747 2805
rect 17494 2796 17500 2848
rect 17552 2796 17558 2848
rect 17604 2836 17632 2876
rect 18800 2836 18828 2944
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 20165 2975 20223 2981
rect 20165 2941 20177 2975
rect 20211 2941 20223 2975
rect 20165 2935 20223 2941
rect 19153 2907 19211 2913
rect 19153 2873 19165 2907
rect 19199 2904 19211 2907
rect 19978 2904 19984 2916
rect 19199 2876 19984 2904
rect 19199 2873 19211 2876
rect 19153 2867 19211 2873
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 17604 2808 18828 2836
rect 19242 2796 19248 2848
rect 19300 2796 19306 2848
rect 1104 2746 24012 2768
rect 1104 2694 1350 2746
rect 1402 2694 1414 2746
rect 1466 2694 1478 2746
rect 1530 2694 1542 2746
rect 1594 2694 1606 2746
rect 1658 2694 4350 2746
rect 4402 2694 4414 2746
rect 4466 2694 4478 2746
rect 4530 2694 4542 2746
rect 4594 2694 4606 2746
rect 4658 2694 7350 2746
rect 7402 2694 7414 2746
rect 7466 2694 7478 2746
rect 7530 2694 7542 2746
rect 7594 2694 7606 2746
rect 7658 2694 10350 2746
rect 10402 2694 10414 2746
rect 10466 2694 10478 2746
rect 10530 2694 10542 2746
rect 10594 2694 10606 2746
rect 10658 2694 13350 2746
rect 13402 2694 13414 2746
rect 13466 2694 13478 2746
rect 13530 2694 13542 2746
rect 13594 2694 13606 2746
rect 13658 2694 16350 2746
rect 16402 2694 16414 2746
rect 16466 2694 16478 2746
rect 16530 2694 16542 2746
rect 16594 2694 16606 2746
rect 16658 2694 19350 2746
rect 19402 2694 19414 2746
rect 19466 2694 19478 2746
rect 19530 2694 19542 2746
rect 19594 2694 19606 2746
rect 19658 2694 22350 2746
rect 22402 2694 22414 2746
rect 22466 2694 22478 2746
rect 22530 2694 22542 2746
rect 22594 2694 22606 2746
rect 22658 2694 24012 2746
rect 1104 2672 24012 2694
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 7190 2632 7196 2644
rect 6135 2604 7196 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 10778 2592 10784 2644
rect 10836 2592 10842 2644
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 12986 2632 12992 2644
rect 11103 2604 12992 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 14424 2604 14473 2632
rect 14424 2592 14430 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15749 2635 15807 2641
rect 15749 2632 15761 2635
rect 15344 2604 15761 2632
rect 15344 2592 15350 2604
rect 15749 2601 15761 2604
rect 15795 2601 15807 2635
rect 15749 2595 15807 2601
rect 16393 2635 16451 2641
rect 16393 2601 16405 2635
rect 16439 2632 16451 2635
rect 16758 2632 16764 2644
rect 16439 2604 16764 2632
rect 16439 2601 16451 2604
rect 16393 2595 16451 2601
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 18322 2632 18328 2644
rect 18187 2604 18328 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 19613 2635 19671 2641
rect 19613 2601 19625 2635
rect 19659 2632 19671 2635
rect 19702 2632 19708 2644
rect 19659 2604 19708 2632
rect 19659 2601 19671 2604
rect 19613 2595 19671 2601
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 8018 2524 8024 2576
rect 8076 2564 8082 2576
rect 11885 2567 11943 2573
rect 8076 2536 9444 2564
rect 8076 2524 8082 2536
rect 8294 2496 8300 2508
rect 7576 2468 8300 2496
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5776 2400 5917 2428
rect 5776 2388 5782 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 6730 2428 6736 2440
rect 6687 2400 6736 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7576 2437 7604 2468
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 9416 2505 9444 2536
rect 11885 2533 11897 2567
rect 11931 2564 11943 2567
rect 12526 2564 12532 2576
rect 11931 2536 12532 2564
rect 11931 2533 11943 2536
rect 11885 2527 11943 2533
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9732 2468 10180 2496
rect 9732 2456 9738 2468
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8628 2400 8677 2428
rect 8628 2388 8634 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9214 2428 9220 2440
rect 9171 2400 9220 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7193 2363 7251 2369
rect 7193 2360 7205 2363
rect 7156 2332 7205 2360
rect 7156 2320 7162 2332
rect 7193 2329 7205 2332
rect 7239 2329 7251 2363
rect 7193 2323 7251 2329
rect 7742 2320 7748 2372
rect 7800 2320 7806 2372
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 10045 2363 10103 2369
rect 10045 2360 10057 2363
rect 9732 2332 10057 2360
rect 9732 2320 9738 2332
rect 10045 2329 10057 2332
rect 10091 2329 10103 2363
rect 10152 2360 10180 2468
rect 17494 2456 17500 2508
rect 17552 2456 17558 2508
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10870 2388 10876 2440
rect 10928 2388 10934 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12802 2428 12808 2440
rect 12759 2400 12808 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14240 2400 14289 2428
rect 14240 2388 14246 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14608 2400 15025 2428
rect 14608 2388 14614 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15528 2400 15577 2428
rect 15528 2388 15534 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16209 2431 16267 2437
rect 16209 2428 16221 2431
rect 16172 2400 16221 2428
rect 16172 2388 16178 2400
rect 16209 2397 16221 2400
rect 16255 2397 16267 2431
rect 16209 2391 16267 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 17512 2428 17540 2456
rect 17267 2400 17540 2428
rect 18325 2431 18383 2437
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 18325 2397 18337 2431
rect 18371 2428 18383 2431
rect 19242 2428 19248 2440
rect 18371 2400 19248 2428
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 21910 2388 21916 2440
rect 21968 2388 21974 2440
rect 10413 2363 10471 2369
rect 10413 2360 10425 2363
rect 10152 2332 10425 2360
rect 10045 2323 10103 2329
rect 10413 2329 10425 2332
rect 10459 2329 10471 2363
rect 10413 2323 10471 2329
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 12308 2332 12357 2360
rect 12308 2320 12314 2332
rect 12345 2329 12357 2332
rect 12391 2329 12403 2363
rect 12345 2323 12403 2329
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 16816 2332 16865 2360
rect 16816 2320 16822 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 16853 2323 16911 2329
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 17497 2363 17555 2369
rect 17497 2360 17509 2363
rect 17460 2332 17509 2360
rect 17460 2320 17466 2332
rect 17497 2329 17509 2332
rect 17543 2329 17555 2363
rect 17497 2323 17555 2329
rect 17865 2363 17923 2369
rect 17865 2329 17877 2363
rect 17911 2360 17923 2363
rect 18414 2360 18420 2372
rect 17911 2332 18420 2360
rect 17911 2329 17923 2332
rect 17865 2323 17923 2329
rect 18414 2320 18420 2332
rect 18472 2320 18478 2372
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14792 2264 15117 2292
rect 14792 2252 14798 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21324 2264 22017 2292
rect 21324 2252 21330 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 1104 2202 24164 2224
rect 1104 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 3042 2202
rect 3094 2150 3106 2202
rect 3158 2150 5850 2202
rect 5902 2150 5914 2202
rect 5966 2150 5978 2202
rect 6030 2150 6042 2202
rect 6094 2150 6106 2202
rect 6158 2150 8850 2202
rect 8902 2150 8914 2202
rect 8966 2150 8978 2202
rect 9030 2150 9042 2202
rect 9094 2150 9106 2202
rect 9158 2150 11850 2202
rect 11902 2150 11914 2202
rect 11966 2150 11978 2202
rect 12030 2150 12042 2202
rect 12094 2150 12106 2202
rect 12158 2150 14850 2202
rect 14902 2150 14914 2202
rect 14966 2150 14978 2202
rect 15030 2150 15042 2202
rect 15094 2150 15106 2202
rect 15158 2150 17850 2202
rect 17902 2150 17914 2202
rect 17966 2150 17978 2202
rect 18030 2150 18042 2202
rect 18094 2150 18106 2202
rect 18158 2150 20850 2202
rect 20902 2150 20914 2202
rect 20966 2150 20978 2202
rect 21030 2150 21042 2202
rect 21094 2150 21106 2202
rect 21158 2150 23850 2202
rect 23902 2150 23914 2202
rect 23966 2150 23978 2202
rect 24030 2150 24042 2202
rect 24094 2150 24106 2202
rect 24158 2150 24164 2202
rect 1104 2128 24164 2150
<< via1 >>
rect 2850 24998 2902 25050
rect 2914 24998 2966 25050
rect 2978 24998 3030 25050
rect 3042 24998 3094 25050
rect 3106 24998 3158 25050
rect 5850 24998 5902 25050
rect 5914 24998 5966 25050
rect 5978 24998 6030 25050
rect 6042 24998 6094 25050
rect 6106 24998 6158 25050
rect 8850 24998 8902 25050
rect 8914 24998 8966 25050
rect 8978 24998 9030 25050
rect 9042 24998 9094 25050
rect 9106 24998 9158 25050
rect 11850 24998 11902 25050
rect 11914 24998 11966 25050
rect 11978 24998 12030 25050
rect 12042 24998 12094 25050
rect 12106 24998 12158 25050
rect 14850 24998 14902 25050
rect 14914 24998 14966 25050
rect 14978 24998 15030 25050
rect 15042 24998 15094 25050
rect 15106 24998 15158 25050
rect 17850 24998 17902 25050
rect 17914 24998 17966 25050
rect 17978 24998 18030 25050
rect 18042 24998 18094 25050
rect 18106 24998 18158 25050
rect 20850 24998 20902 25050
rect 20914 24998 20966 25050
rect 20978 24998 21030 25050
rect 21042 24998 21094 25050
rect 21106 24998 21158 25050
rect 23850 24998 23902 25050
rect 23914 24998 23966 25050
rect 23978 24998 24030 25050
rect 24042 24998 24094 25050
rect 24106 24998 24158 25050
rect 9312 24828 9364 24880
rect 5172 24760 5224 24812
rect 5632 24735 5684 24744
rect 5632 24701 5641 24735
rect 5641 24701 5675 24735
rect 5675 24701 5684 24735
rect 5632 24692 5684 24701
rect 6552 24692 6604 24744
rect 7196 24760 7248 24812
rect 8392 24760 8444 24812
rect 7840 24692 7892 24744
rect 9680 24760 9732 24812
rect 10140 24692 10192 24744
rect 5172 24624 5224 24676
rect 5724 24624 5776 24676
rect 10324 24624 10376 24676
rect 12440 24760 12492 24812
rect 12900 24760 12952 24812
rect 10784 24735 10836 24744
rect 10784 24701 10793 24735
rect 10793 24701 10827 24735
rect 10827 24701 10836 24735
rect 10784 24692 10836 24701
rect 11428 24692 11480 24744
rect 12256 24692 12308 24744
rect 13544 24760 13596 24812
rect 14740 24760 14792 24812
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 15476 24760 15528 24812
rect 16212 24760 16264 24812
rect 14648 24735 14700 24744
rect 14648 24701 14657 24735
rect 14657 24701 14691 24735
rect 14691 24701 14700 24735
rect 14648 24692 14700 24701
rect 16028 24692 16080 24744
rect 18788 24760 18840 24812
rect 19340 24760 19392 24812
rect 19064 24692 19116 24744
rect 19248 24692 19300 24744
rect 19984 24760 20036 24812
rect 20444 24803 20496 24812
rect 20444 24769 20453 24803
rect 20453 24769 20487 24803
rect 20487 24769 20496 24803
rect 20444 24760 20496 24769
rect 11520 24624 11572 24676
rect 12900 24624 12952 24676
rect 4988 24599 5040 24608
rect 4988 24565 4997 24599
rect 4997 24565 5031 24599
rect 5031 24565 5040 24599
rect 4988 24556 5040 24565
rect 6460 24556 6512 24608
rect 7104 24556 7156 24608
rect 8668 24556 8720 24608
rect 9312 24599 9364 24608
rect 9312 24565 9321 24599
rect 9321 24565 9355 24599
rect 9355 24565 9364 24599
rect 9312 24556 9364 24565
rect 9404 24599 9456 24608
rect 9404 24565 9413 24599
rect 9413 24565 9447 24599
rect 9447 24565 9456 24599
rect 9404 24556 9456 24565
rect 9496 24556 9548 24608
rect 11612 24556 11664 24608
rect 13268 24556 13320 24608
rect 13820 24599 13872 24608
rect 13820 24565 13829 24599
rect 13829 24565 13863 24599
rect 13863 24565 13872 24599
rect 13820 24556 13872 24565
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 16120 24556 16172 24608
rect 18328 24556 18380 24608
rect 18972 24556 19024 24608
rect 19156 24556 19208 24608
rect 20720 24556 20772 24608
rect 1350 24454 1402 24506
rect 1414 24454 1466 24506
rect 1478 24454 1530 24506
rect 1542 24454 1594 24506
rect 1606 24454 1658 24506
rect 4350 24454 4402 24506
rect 4414 24454 4466 24506
rect 4478 24454 4530 24506
rect 4542 24454 4594 24506
rect 4606 24454 4658 24506
rect 7350 24454 7402 24506
rect 7414 24454 7466 24506
rect 7478 24454 7530 24506
rect 7542 24454 7594 24506
rect 7606 24454 7658 24506
rect 10350 24454 10402 24506
rect 10414 24454 10466 24506
rect 10478 24454 10530 24506
rect 10542 24454 10594 24506
rect 10606 24454 10658 24506
rect 13350 24454 13402 24506
rect 13414 24454 13466 24506
rect 13478 24454 13530 24506
rect 13542 24454 13594 24506
rect 13606 24454 13658 24506
rect 16350 24454 16402 24506
rect 16414 24454 16466 24506
rect 16478 24454 16530 24506
rect 16542 24454 16594 24506
rect 16606 24454 16658 24506
rect 19350 24454 19402 24506
rect 19414 24454 19466 24506
rect 19478 24454 19530 24506
rect 19542 24454 19594 24506
rect 19606 24454 19658 24506
rect 22350 24454 22402 24506
rect 22414 24454 22466 24506
rect 22478 24454 22530 24506
rect 22542 24454 22594 24506
rect 22606 24454 22658 24506
rect 6736 24352 6788 24404
rect 10968 24352 11020 24404
rect 12440 24395 12492 24404
rect 12440 24361 12449 24395
rect 12449 24361 12483 24395
rect 12483 24361 12492 24395
rect 12440 24352 12492 24361
rect 16212 24395 16264 24404
rect 16212 24361 16221 24395
rect 16221 24361 16255 24395
rect 16255 24361 16264 24395
rect 16212 24352 16264 24361
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 5632 24284 5684 24336
rect 19064 24284 19116 24336
rect 9220 24216 9272 24268
rect 13728 24259 13780 24268
rect 13728 24225 13737 24259
rect 13737 24225 13771 24259
rect 13771 24225 13780 24259
rect 13728 24216 13780 24225
rect 16212 24216 16264 24268
rect 18236 24216 18288 24268
rect 19156 24216 19208 24268
rect 3516 24148 3568 24200
rect 3424 24080 3476 24132
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 5448 24012 5500 24064
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 7932 24080 7984 24132
rect 8760 24148 8812 24200
rect 9312 24148 9364 24200
rect 7012 24055 7064 24064
rect 7012 24021 7021 24055
rect 7021 24021 7055 24055
rect 7055 24021 7064 24055
rect 7012 24012 7064 24021
rect 7288 24055 7340 24064
rect 7288 24021 7297 24055
rect 7297 24021 7331 24055
rect 7331 24021 7340 24055
rect 7288 24012 7340 24021
rect 8392 24012 8444 24064
rect 8760 24055 8812 24064
rect 8760 24021 8769 24055
rect 8769 24021 8803 24055
rect 8803 24021 8812 24055
rect 8760 24012 8812 24021
rect 9312 24055 9364 24064
rect 9312 24021 9321 24055
rect 9321 24021 9355 24055
rect 9355 24021 9364 24055
rect 9312 24012 9364 24021
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 9864 24080 9916 24132
rect 11704 24080 11756 24132
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 13084 24080 13136 24132
rect 9588 24012 9640 24064
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 12532 24012 12584 24064
rect 12716 24055 12768 24064
rect 12716 24021 12725 24055
rect 12725 24021 12759 24055
rect 12759 24021 12768 24055
rect 12716 24012 12768 24021
rect 14096 24148 14148 24200
rect 14188 24191 14240 24200
rect 14188 24157 14197 24191
rect 14197 24157 14231 24191
rect 14231 24157 14240 24191
rect 14188 24148 14240 24157
rect 14280 24148 14332 24200
rect 13912 24080 13964 24132
rect 16580 24080 16632 24132
rect 16856 24080 16908 24132
rect 18420 24080 18472 24132
rect 18972 24080 19024 24132
rect 19616 24080 19668 24132
rect 20168 24080 20220 24132
rect 20260 24080 20312 24132
rect 13820 24012 13872 24064
rect 14372 24055 14424 24064
rect 14372 24021 14381 24055
rect 14381 24021 14415 24055
rect 14415 24021 14424 24055
rect 14372 24012 14424 24021
rect 14556 24012 14608 24064
rect 15568 24012 15620 24064
rect 18880 24012 18932 24064
rect 2850 23910 2902 23962
rect 2914 23910 2966 23962
rect 2978 23910 3030 23962
rect 3042 23910 3094 23962
rect 3106 23910 3158 23962
rect 5850 23910 5902 23962
rect 5914 23910 5966 23962
rect 5978 23910 6030 23962
rect 6042 23910 6094 23962
rect 6106 23910 6158 23962
rect 8850 23910 8902 23962
rect 8914 23910 8966 23962
rect 8978 23910 9030 23962
rect 9042 23910 9094 23962
rect 9106 23910 9158 23962
rect 11850 23910 11902 23962
rect 11914 23910 11966 23962
rect 11978 23910 12030 23962
rect 12042 23910 12094 23962
rect 12106 23910 12158 23962
rect 14850 23910 14902 23962
rect 14914 23910 14966 23962
rect 14978 23910 15030 23962
rect 15042 23910 15094 23962
rect 15106 23910 15158 23962
rect 17850 23910 17902 23962
rect 17914 23910 17966 23962
rect 17978 23910 18030 23962
rect 18042 23910 18094 23962
rect 18106 23910 18158 23962
rect 20850 23910 20902 23962
rect 20914 23910 20966 23962
rect 20978 23910 21030 23962
rect 21042 23910 21094 23962
rect 21106 23910 21158 23962
rect 23850 23910 23902 23962
rect 23914 23910 23966 23962
rect 23978 23910 24030 23962
rect 24042 23910 24094 23962
rect 24106 23910 24158 23962
rect 3424 23851 3476 23860
rect 3424 23817 3433 23851
rect 3433 23817 3467 23851
rect 3467 23817 3476 23851
rect 3424 23808 3476 23817
rect 5448 23808 5500 23860
rect 5724 23851 5776 23860
rect 5724 23817 5733 23851
rect 5733 23817 5767 23851
rect 5767 23817 5776 23851
rect 5724 23808 5776 23817
rect 7104 23808 7156 23860
rect 4252 23740 4304 23792
rect 7288 23740 7340 23792
rect 8300 23740 8352 23792
rect 9864 23851 9916 23860
rect 9864 23817 9873 23851
rect 9873 23817 9907 23851
rect 9907 23817 9916 23851
rect 9864 23808 9916 23817
rect 11428 23808 11480 23860
rect 14648 23808 14700 23860
rect 15844 23808 15896 23860
rect 16580 23808 16632 23860
rect 12716 23740 12768 23792
rect 13912 23783 13964 23792
rect 13912 23749 13921 23783
rect 13921 23749 13955 23783
rect 13955 23749 13964 23783
rect 13912 23740 13964 23749
rect 19616 23740 19668 23792
rect 20444 23808 20496 23860
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 3792 23715 3844 23724
rect 3792 23681 3826 23715
rect 3826 23681 3844 23715
rect 3792 23672 3844 23681
rect 6736 23672 6788 23724
rect 9496 23672 9548 23724
rect 9680 23715 9732 23724
rect 9680 23681 9689 23715
rect 9689 23681 9723 23715
rect 9723 23681 9732 23715
rect 9680 23672 9732 23681
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 6276 23604 6328 23656
rect 7932 23647 7984 23656
rect 7932 23613 7941 23647
rect 7941 23613 7975 23647
rect 7975 23613 7984 23647
rect 7932 23604 7984 23613
rect 10784 23672 10836 23724
rect 11336 23672 11388 23724
rect 11888 23672 11940 23724
rect 5632 23468 5684 23520
rect 6092 23468 6144 23520
rect 6552 23536 6604 23588
rect 6460 23468 6512 23520
rect 12256 23647 12308 23656
rect 12256 23613 12265 23647
rect 12265 23613 12299 23647
rect 12299 23613 12308 23647
rect 12256 23604 12308 23613
rect 14648 23672 14700 23724
rect 14832 23715 14884 23724
rect 14832 23681 14841 23715
rect 14841 23681 14875 23715
rect 14875 23681 14884 23715
rect 14832 23672 14884 23681
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 16764 23672 16816 23724
rect 10140 23468 10192 23520
rect 10876 23468 10928 23520
rect 11520 23511 11572 23520
rect 11520 23477 11529 23511
rect 11529 23477 11563 23511
rect 11563 23477 11572 23511
rect 11520 23468 11572 23477
rect 15752 23647 15804 23656
rect 15752 23613 15761 23647
rect 15761 23613 15795 23647
rect 15795 23613 15804 23647
rect 15752 23604 15804 23613
rect 17592 23647 17644 23656
rect 17592 23613 17601 23647
rect 17601 23613 17635 23647
rect 17635 23613 17644 23647
rect 17592 23604 17644 23613
rect 17684 23647 17736 23656
rect 17684 23613 17693 23647
rect 17693 23613 17727 23647
rect 17727 23613 17736 23647
rect 17684 23604 17736 23613
rect 18420 23604 18472 23656
rect 18604 23647 18656 23656
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 18696 23604 18748 23656
rect 19064 23604 19116 23656
rect 19248 23604 19300 23656
rect 19984 23604 20036 23656
rect 20444 23647 20496 23656
rect 20444 23613 20453 23647
rect 20453 23613 20487 23647
rect 20487 23613 20496 23647
rect 20444 23604 20496 23613
rect 15108 23579 15160 23588
rect 15108 23545 15117 23579
rect 15117 23545 15151 23579
rect 15151 23545 15160 23579
rect 15108 23536 15160 23545
rect 15476 23468 15528 23520
rect 17316 23468 17368 23520
rect 19156 23579 19208 23588
rect 19156 23545 19165 23579
rect 19165 23545 19199 23579
rect 19199 23545 19208 23579
rect 19156 23536 19208 23545
rect 18604 23468 18656 23520
rect 19892 23511 19944 23520
rect 19892 23477 19901 23511
rect 19901 23477 19935 23511
rect 19935 23477 19944 23511
rect 19892 23468 19944 23477
rect 1350 23366 1402 23418
rect 1414 23366 1466 23418
rect 1478 23366 1530 23418
rect 1542 23366 1594 23418
rect 1606 23366 1658 23418
rect 4350 23366 4402 23418
rect 4414 23366 4466 23418
rect 4478 23366 4530 23418
rect 4542 23366 4594 23418
rect 4606 23366 4658 23418
rect 7350 23366 7402 23418
rect 7414 23366 7466 23418
rect 7478 23366 7530 23418
rect 7542 23366 7594 23418
rect 7606 23366 7658 23418
rect 10350 23366 10402 23418
rect 10414 23366 10466 23418
rect 10478 23366 10530 23418
rect 10542 23366 10594 23418
rect 10606 23366 10658 23418
rect 13350 23366 13402 23418
rect 13414 23366 13466 23418
rect 13478 23366 13530 23418
rect 13542 23366 13594 23418
rect 13606 23366 13658 23418
rect 16350 23366 16402 23418
rect 16414 23366 16466 23418
rect 16478 23366 16530 23418
rect 16542 23366 16594 23418
rect 16606 23366 16658 23418
rect 19350 23366 19402 23418
rect 19414 23366 19466 23418
rect 19478 23366 19530 23418
rect 19542 23366 19594 23418
rect 19606 23366 19658 23418
rect 22350 23366 22402 23418
rect 22414 23366 22466 23418
rect 22478 23366 22530 23418
rect 22542 23366 22594 23418
rect 22606 23366 22658 23418
rect 3792 23264 3844 23316
rect 6552 23196 6604 23248
rect 5264 23128 5316 23180
rect 5448 23128 5500 23180
rect 5908 23128 5960 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 6644 23128 6696 23180
rect 7840 23239 7892 23248
rect 7840 23205 7849 23239
rect 7849 23205 7883 23239
rect 7883 23205 7892 23239
rect 7840 23196 7892 23205
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 12164 23264 12216 23316
rect 14740 23264 14792 23316
rect 15660 23264 15712 23316
rect 16764 23264 16816 23316
rect 18696 23264 18748 23316
rect 11244 23239 11296 23248
rect 11244 23205 11253 23239
rect 11253 23205 11287 23239
rect 11287 23205 11296 23239
rect 11244 23196 11296 23205
rect 11428 23196 11480 23248
rect 9404 23171 9456 23180
rect 9404 23137 9413 23171
rect 9413 23137 9447 23171
rect 9447 23137 9456 23171
rect 9404 23128 9456 23137
rect 9496 23171 9548 23180
rect 9496 23137 9505 23171
rect 9505 23137 9539 23171
rect 9539 23137 9548 23171
rect 9496 23128 9548 23137
rect 10048 23128 10100 23180
rect 11888 23171 11940 23180
rect 11888 23137 11897 23171
rect 11897 23137 11931 23171
rect 11931 23137 11940 23171
rect 11888 23128 11940 23137
rect 15568 23128 15620 23180
rect 15844 23171 15896 23180
rect 15844 23137 15853 23171
rect 15853 23137 15887 23171
rect 15887 23137 15896 23171
rect 15844 23128 15896 23137
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 10876 23103 10928 23112
rect 10876 23069 10894 23103
rect 10894 23069 10928 23103
rect 10876 23060 10928 23069
rect 4712 22967 4764 22976
rect 4712 22933 4721 22967
rect 4721 22933 4755 22967
rect 4755 22933 4764 22967
rect 4712 22924 4764 22933
rect 4804 22967 4856 22976
rect 4804 22933 4813 22967
rect 4813 22933 4847 22967
rect 4847 22933 4856 22967
rect 4804 22924 4856 22933
rect 6644 22924 6696 22976
rect 6828 22924 6880 22976
rect 9496 22924 9548 22976
rect 9956 22924 10008 22976
rect 12256 23060 12308 23112
rect 12440 23103 12492 23112
rect 12440 23069 12474 23103
rect 12474 23069 12492 23103
rect 12440 23060 12492 23069
rect 15200 23060 15252 23112
rect 16212 23060 16264 23112
rect 18420 23171 18472 23180
rect 18420 23137 18429 23171
rect 18429 23137 18463 23171
rect 18463 23137 18472 23171
rect 18420 23128 18472 23137
rect 18512 23171 18564 23180
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 18236 23060 18288 23112
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 19892 23264 19944 23316
rect 19984 23264 20036 23316
rect 18972 23060 19024 23112
rect 14372 23035 14424 23044
rect 14372 23001 14406 23035
rect 14406 23001 14424 23035
rect 14372 22992 14424 23001
rect 14648 22992 14700 23044
rect 17132 22992 17184 23044
rect 17224 22992 17276 23044
rect 15752 22924 15804 22976
rect 16396 22924 16448 22976
rect 2850 22822 2902 22874
rect 2914 22822 2966 22874
rect 2978 22822 3030 22874
rect 3042 22822 3094 22874
rect 3106 22822 3158 22874
rect 5850 22822 5902 22874
rect 5914 22822 5966 22874
rect 5978 22822 6030 22874
rect 6042 22822 6094 22874
rect 6106 22822 6158 22874
rect 8850 22822 8902 22874
rect 8914 22822 8966 22874
rect 8978 22822 9030 22874
rect 9042 22822 9094 22874
rect 9106 22822 9158 22874
rect 11850 22822 11902 22874
rect 11914 22822 11966 22874
rect 11978 22822 12030 22874
rect 12042 22822 12094 22874
rect 12106 22822 12158 22874
rect 14850 22822 14902 22874
rect 14914 22822 14966 22874
rect 14978 22822 15030 22874
rect 15042 22822 15094 22874
rect 15106 22822 15158 22874
rect 17850 22822 17902 22874
rect 17914 22822 17966 22874
rect 17978 22822 18030 22874
rect 18042 22822 18094 22874
rect 18106 22822 18158 22874
rect 20850 22822 20902 22874
rect 20914 22822 20966 22874
rect 20978 22822 21030 22874
rect 21042 22822 21094 22874
rect 21106 22822 21158 22874
rect 23850 22822 23902 22874
rect 23914 22822 23966 22874
rect 23978 22822 24030 22874
rect 24042 22822 24094 22874
rect 24106 22822 24158 22874
rect 4252 22763 4304 22772
rect 4252 22729 4261 22763
rect 4261 22729 4295 22763
rect 4295 22729 4304 22763
rect 4252 22720 4304 22729
rect 4712 22720 4764 22772
rect 6276 22720 6328 22772
rect 6736 22763 6788 22772
rect 6736 22729 6745 22763
rect 6745 22729 6779 22763
rect 6779 22729 6788 22763
rect 6736 22720 6788 22729
rect 6828 22763 6880 22772
rect 6828 22729 6837 22763
rect 6837 22729 6871 22763
rect 6871 22729 6880 22763
rect 6828 22720 6880 22729
rect 9312 22720 9364 22772
rect 9680 22720 9732 22772
rect 11520 22720 11572 22772
rect 13084 22763 13136 22772
rect 13084 22729 13093 22763
rect 13093 22729 13127 22763
rect 13127 22729 13136 22763
rect 13084 22720 13136 22729
rect 14188 22720 14240 22772
rect 14648 22763 14700 22772
rect 14648 22729 14657 22763
rect 14657 22729 14691 22763
rect 14691 22729 14700 22763
rect 14648 22720 14700 22729
rect 16856 22763 16908 22772
rect 16856 22729 16865 22763
rect 16865 22729 16899 22763
rect 16899 22729 16908 22763
rect 16856 22720 16908 22729
rect 17132 22763 17184 22772
rect 17132 22729 17141 22763
rect 17141 22729 17175 22763
rect 17175 22729 17184 22763
rect 17132 22720 17184 22729
rect 17592 22720 17644 22772
rect 20260 22720 20312 22772
rect 4804 22652 4856 22704
rect 5264 22652 5316 22704
rect 4988 22584 5040 22636
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 6368 22584 6420 22636
rect 8392 22652 8444 22704
rect 9496 22652 9548 22704
rect 9220 22584 9272 22636
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 13820 22584 13872 22636
rect 14648 22584 14700 22636
rect 17224 22584 17276 22636
rect 17316 22627 17368 22636
rect 17316 22593 17325 22627
rect 17325 22593 17359 22627
rect 17359 22593 17368 22627
rect 17316 22584 17368 22593
rect 18696 22584 18748 22636
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 4896 22559 4948 22568
rect 4896 22525 4905 22559
rect 4905 22525 4939 22559
rect 4939 22525 4948 22559
rect 4896 22516 4948 22525
rect 6828 22516 6880 22568
rect 7932 22559 7984 22568
rect 7932 22525 7941 22559
rect 7941 22525 7975 22559
rect 7975 22525 7984 22559
rect 7932 22516 7984 22525
rect 5080 22380 5132 22432
rect 14372 22516 14424 22568
rect 15660 22559 15712 22568
rect 15660 22525 15669 22559
rect 15669 22525 15703 22559
rect 15703 22525 15712 22559
rect 15660 22516 15712 22525
rect 16396 22559 16448 22568
rect 16396 22525 16405 22559
rect 16405 22525 16439 22559
rect 16439 22525 16448 22559
rect 16396 22516 16448 22525
rect 14280 22380 14332 22432
rect 14648 22380 14700 22432
rect 1350 22278 1402 22330
rect 1414 22278 1466 22330
rect 1478 22278 1530 22330
rect 1542 22278 1594 22330
rect 1606 22278 1658 22330
rect 4350 22278 4402 22330
rect 4414 22278 4466 22330
rect 4478 22278 4530 22330
rect 4542 22278 4594 22330
rect 4606 22278 4658 22330
rect 7350 22278 7402 22330
rect 7414 22278 7466 22330
rect 7478 22278 7530 22330
rect 7542 22278 7594 22330
rect 7606 22278 7658 22330
rect 10350 22278 10402 22330
rect 10414 22278 10466 22330
rect 10478 22278 10530 22330
rect 10542 22278 10594 22330
rect 10606 22278 10658 22330
rect 13350 22278 13402 22330
rect 13414 22278 13466 22330
rect 13478 22278 13530 22330
rect 13542 22278 13594 22330
rect 13606 22278 13658 22330
rect 16350 22278 16402 22330
rect 16414 22278 16466 22330
rect 16478 22278 16530 22330
rect 16542 22278 16594 22330
rect 16606 22278 16658 22330
rect 19350 22278 19402 22330
rect 19414 22278 19466 22330
rect 19478 22278 19530 22330
rect 19542 22278 19594 22330
rect 19606 22278 19658 22330
rect 22350 22278 22402 22330
rect 22414 22278 22466 22330
rect 22478 22278 22530 22330
rect 22542 22278 22594 22330
rect 22606 22278 22658 22330
rect 4896 22176 4948 22228
rect 5172 22040 5224 22092
rect 9404 22176 9456 22228
rect 9220 22108 9272 22160
rect 4620 22015 4672 22024
rect 4620 21981 4629 22015
rect 4629 21981 4663 22015
rect 4663 21981 4672 22015
rect 4620 21972 4672 21981
rect 4804 21904 4856 21956
rect 5632 21972 5684 22024
rect 7932 22040 7984 22092
rect 13728 22108 13780 22160
rect 18420 22108 18472 22160
rect 14188 22040 14240 22092
rect 14372 22040 14424 22092
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 8760 21972 8812 22024
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 11520 21972 11572 22024
rect 6736 21904 6788 21956
rect 7656 21947 7708 21956
rect 7656 21913 7665 21947
rect 7665 21913 7699 21947
rect 7699 21913 7708 21947
rect 7656 21904 7708 21913
rect 13176 21972 13228 22024
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 15384 21972 15436 21981
rect 16672 22015 16724 22024
rect 16672 21981 16681 22015
rect 16681 21981 16715 22015
rect 16715 21981 16724 22015
rect 16672 21972 16724 21981
rect 19248 21972 19300 22024
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 14004 21904 14056 21956
rect 16304 21904 16356 21956
rect 18972 21904 19024 21956
rect 4252 21836 4304 21888
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 8024 21836 8076 21888
rect 9220 21836 9272 21888
rect 10232 21836 10284 21888
rect 12532 21836 12584 21888
rect 12716 21879 12768 21888
rect 12716 21845 12725 21879
rect 12725 21845 12759 21879
rect 12759 21845 12768 21879
rect 12716 21836 12768 21845
rect 13544 21836 13596 21888
rect 14464 21836 14516 21888
rect 15660 21836 15712 21888
rect 18512 21836 18564 21888
rect 18604 21836 18656 21888
rect 2850 21734 2902 21786
rect 2914 21734 2966 21786
rect 2978 21734 3030 21786
rect 3042 21734 3094 21786
rect 3106 21734 3158 21786
rect 5850 21734 5902 21786
rect 5914 21734 5966 21786
rect 5978 21734 6030 21786
rect 6042 21734 6094 21786
rect 6106 21734 6158 21786
rect 8850 21734 8902 21786
rect 8914 21734 8966 21786
rect 8978 21734 9030 21786
rect 9042 21734 9094 21786
rect 9106 21734 9158 21786
rect 11850 21734 11902 21786
rect 11914 21734 11966 21786
rect 11978 21734 12030 21786
rect 12042 21734 12094 21786
rect 12106 21734 12158 21786
rect 14850 21734 14902 21786
rect 14914 21734 14966 21786
rect 14978 21734 15030 21786
rect 15042 21734 15094 21786
rect 15106 21734 15158 21786
rect 17850 21734 17902 21786
rect 17914 21734 17966 21786
rect 17978 21734 18030 21786
rect 18042 21734 18094 21786
rect 18106 21734 18158 21786
rect 20850 21734 20902 21786
rect 20914 21734 20966 21786
rect 20978 21734 21030 21786
rect 21042 21734 21094 21786
rect 21106 21734 21158 21786
rect 23850 21734 23902 21786
rect 23914 21734 23966 21786
rect 23978 21734 24030 21786
rect 24042 21734 24094 21786
rect 24106 21734 24158 21786
rect 6368 21675 6420 21684
rect 6368 21641 6377 21675
rect 6377 21641 6411 21675
rect 6411 21641 6420 21675
rect 6368 21632 6420 21641
rect 11520 21675 11572 21684
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 13176 21675 13228 21684
rect 13176 21641 13185 21675
rect 13185 21641 13219 21675
rect 13219 21641 13228 21675
rect 13176 21632 13228 21641
rect 13544 21675 13596 21684
rect 13544 21641 13553 21675
rect 13553 21641 13587 21675
rect 13587 21641 13596 21675
rect 13544 21632 13596 21641
rect 14004 21675 14056 21684
rect 14004 21641 14013 21675
rect 14013 21641 14047 21675
rect 14047 21641 14056 21675
rect 14004 21632 14056 21641
rect 14464 21675 14516 21684
rect 14464 21641 14473 21675
rect 14473 21641 14507 21675
rect 14507 21641 14516 21675
rect 14464 21632 14516 21641
rect 14648 21632 14700 21684
rect 16672 21632 16724 21684
rect 5172 21607 5224 21616
rect 5172 21573 5181 21607
rect 5181 21573 5215 21607
rect 5215 21573 5224 21607
rect 5172 21564 5224 21573
rect 9404 21564 9456 21616
rect 17684 21632 17736 21684
rect 18604 21675 18656 21684
rect 18604 21641 18613 21675
rect 18613 21641 18647 21675
rect 18647 21641 18656 21675
rect 18604 21632 18656 21641
rect 18696 21632 18748 21684
rect 20444 21632 20496 21684
rect 3792 21496 3844 21548
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 8852 21496 8904 21548
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 5448 21428 5500 21480
rect 6644 21428 6696 21480
rect 7012 21428 7064 21480
rect 7932 21428 7984 21480
rect 9680 21428 9732 21480
rect 14464 21496 14516 21548
rect 11520 21428 11572 21480
rect 11428 21360 11480 21412
rect 13728 21471 13780 21480
rect 13728 21437 13737 21471
rect 13737 21437 13771 21471
rect 13771 21437 13780 21471
rect 13728 21428 13780 21437
rect 14188 21428 14240 21480
rect 16120 21539 16172 21548
rect 16120 21505 16138 21539
rect 16138 21505 16172 21539
rect 16120 21496 16172 21505
rect 16304 21496 16356 21548
rect 16856 21496 16908 21548
rect 18788 21496 18840 21548
rect 18972 21496 19024 21548
rect 19248 21496 19300 21548
rect 19984 21496 20036 21548
rect 21272 21496 21324 21548
rect 4160 21292 4212 21344
rect 4620 21335 4672 21344
rect 4620 21301 4629 21335
rect 4629 21301 4663 21335
rect 4663 21301 4672 21335
rect 4620 21292 4672 21301
rect 6092 21292 6144 21344
rect 10140 21292 10192 21344
rect 10324 21292 10376 21344
rect 11336 21335 11388 21344
rect 11336 21301 11345 21335
rect 11345 21301 11379 21335
rect 11379 21301 11388 21335
rect 11336 21292 11388 21301
rect 14556 21292 14608 21344
rect 18604 21428 18656 21480
rect 19156 21292 19208 21344
rect 19800 21292 19852 21344
rect 21180 21292 21232 21344
rect 23572 21335 23624 21344
rect 23572 21301 23581 21335
rect 23581 21301 23615 21335
rect 23615 21301 23624 21335
rect 23572 21292 23624 21301
rect 1350 21190 1402 21242
rect 1414 21190 1466 21242
rect 1478 21190 1530 21242
rect 1542 21190 1594 21242
rect 1606 21190 1658 21242
rect 4350 21190 4402 21242
rect 4414 21190 4466 21242
rect 4478 21190 4530 21242
rect 4542 21190 4594 21242
rect 4606 21190 4658 21242
rect 7350 21190 7402 21242
rect 7414 21190 7466 21242
rect 7478 21190 7530 21242
rect 7542 21190 7594 21242
rect 7606 21190 7658 21242
rect 10350 21190 10402 21242
rect 10414 21190 10466 21242
rect 10478 21190 10530 21242
rect 10542 21190 10594 21242
rect 10606 21190 10658 21242
rect 13350 21190 13402 21242
rect 13414 21190 13466 21242
rect 13478 21190 13530 21242
rect 13542 21190 13594 21242
rect 13606 21190 13658 21242
rect 16350 21190 16402 21242
rect 16414 21190 16466 21242
rect 16478 21190 16530 21242
rect 16542 21190 16594 21242
rect 16606 21190 16658 21242
rect 19350 21190 19402 21242
rect 19414 21190 19466 21242
rect 19478 21190 19530 21242
rect 19542 21190 19594 21242
rect 19606 21190 19658 21242
rect 22350 21190 22402 21242
rect 22414 21190 22466 21242
rect 22478 21190 22530 21242
rect 22542 21190 22594 21242
rect 22606 21190 22658 21242
rect 3792 21131 3844 21140
rect 3792 21097 3801 21131
rect 3801 21097 3835 21131
rect 3835 21097 3844 21131
rect 3792 21088 3844 21097
rect 4712 21088 4764 21140
rect 8852 21088 8904 21140
rect 10140 21088 10192 21140
rect 6552 21020 6604 21072
rect 5264 20952 5316 21004
rect 5632 20952 5684 21004
rect 6092 20995 6144 21004
rect 6092 20961 6101 20995
rect 6101 20961 6135 20995
rect 6135 20961 6144 20995
rect 6092 20952 6144 20961
rect 6276 20952 6328 21004
rect 7012 20995 7064 21004
rect 7012 20961 7021 20995
rect 7021 20961 7055 20995
rect 7055 20961 7064 20995
rect 7012 20952 7064 20961
rect 9312 20952 9364 21004
rect 14096 21088 14148 21140
rect 13636 21063 13688 21072
rect 13636 21029 13645 21063
rect 13645 21029 13679 21063
rect 13679 21029 13688 21063
rect 13636 21020 13688 21029
rect 3516 20748 3568 20800
rect 4252 20884 4304 20936
rect 4804 20884 4856 20936
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6644 20748 6696 20800
rect 7932 20884 7984 20936
rect 8760 20927 8812 20936
rect 8760 20893 8769 20927
rect 8769 20893 8803 20927
rect 8803 20893 8812 20927
rect 8760 20884 8812 20893
rect 9220 20884 9272 20936
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10876 20952 10928 21004
rect 11336 20952 11388 21004
rect 14556 21020 14608 21072
rect 15108 21088 15160 21140
rect 15384 21088 15436 21140
rect 16028 21088 16080 21140
rect 16856 21088 16908 21140
rect 20352 21088 20404 21140
rect 18972 21020 19024 21072
rect 15108 20995 15160 21004
rect 15108 20961 15142 20995
rect 15142 20961 15160 20995
rect 15108 20952 15160 20961
rect 15476 20952 15528 21004
rect 15844 20952 15896 21004
rect 18420 20952 18472 21004
rect 19064 20952 19116 21004
rect 21180 20995 21232 21004
rect 21180 20961 21189 20995
rect 21189 20961 21223 20995
rect 21223 20961 21232 20995
rect 21180 20952 21232 20961
rect 21364 20995 21416 21004
rect 21364 20961 21373 20995
rect 21373 20961 21407 20995
rect 21407 20961 21416 20995
rect 21364 20952 21416 20961
rect 8024 20816 8076 20868
rect 11244 20927 11296 20936
rect 11244 20893 11253 20927
rect 11253 20893 11287 20927
rect 11287 20893 11296 20927
rect 11244 20884 11296 20893
rect 11428 20816 11480 20868
rect 12532 20927 12584 20936
rect 12532 20893 12566 20927
rect 12566 20893 12584 20927
rect 12532 20884 12584 20893
rect 13912 20884 13964 20936
rect 7104 20791 7156 20800
rect 7104 20757 7113 20791
rect 7113 20757 7147 20791
rect 7147 20757 7156 20791
rect 7104 20748 7156 20757
rect 8576 20791 8628 20800
rect 8576 20757 8585 20791
rect 8585 20757 8619 20791
rect 8619 20757 8628 20791
rect 8576 20748 8628 20757
rect 11152 20748 11204 20800
rect 11244 20748 11296 20800
rect 14004 20748 14056 20800
rect 15016 20927 15068 20936
rect 15016 20893 15025 20927
rect 15025 20893 15059 20927
rect 15059 20893 15068 20927
rect 15016 20884 15068 20893
rect 16488 20884 16540 20936
rect 16948 20859 17000 20868
rect 16948 20825 16982 20859
rect 16982 20825 17000 20859
rect 16948 20816 17000 20825
rect 15384 20748 15436 20800
rect 18512 20927 18564 20936
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 20720 20884 20772 20936
rect 19708 20816 19760 20868
rect 18604 20791 18656 20800
rect 18604 20757 18613 20791
rect 18613 20757 18647 20791
rect 18647 20757 18656 20791
rect 18604 20748 18656 20757
rect 20720 20791 20772 20800
rect 20720 20757 20729 20791
rect 20729 20757 20763 20791
rect 20763 20757 20772 20791
rect 20720 20748 20772 20757
rect 2850 20646 2902 20698
rect 2914 20646 2966 20698
rect 2978 20646 3030 20698
rect 3042 20646 3094 20698
rect 3106 20646 3158 20698
rect 5850 20646 5902 20698
rect 5914 20646 5966 20698
rect 5978 20646 6030 20698
rect 6042 20646 6094 20698
rect 6106 20646 6158 20698
rect 8850 20646 8902 20698
rect 8914 20646 8966 20698
rect 8978 20646 9030 20698
rect 9042 20646 9094 20698
rect 9106 20646 9158 20698
rect 11850 20646 11902 20698
rect 11914 20646 11966 20698
rect 11978 20646 12030 20698
rect 12042 20646 12094 20698
rect 12106 20646 12158 20698
rect 14850 20646 14902 20698
rect 14914 20646 14966 20698
rect 14978 20646 15030 20698
rect 15042 20646 15094 20698
rect 15106 20646 15158 20698
rect 17850 20646 17902 20698
rect 17914 20646 17966 20698
rect 17978 20646 18030 20698
rect 18042 20646 18094 20698
rect 18106 20646 18158 20698
rect 20850 20646 20902 20698
rect 20914 20646 20966 20698
rect 20978 20646 21030 20698
rect 21042 20646 21094 20698
rect 21106 20646 21158 20698
rect 23850 20646 23902 20698
rect 23914 20646 23966 20698
rect 23978 20646 24030 20698
rect 24042 20646 24094 20698
rect 24106 20646 24158 20698
rect 5632 20544 5684 20596
rect 7012 20544 7064 20596
rect 7748 20544 7800 20596
rect 9312 20587 9364 20596
rect 9312 20553 9321 20587
rect 9321 20553 9355 20587
rect 9355 20553 9364 20587
rect 9312 20544 9364 20553
rect 3516 20451 3568 20460
rect 3516 20417 3550 20451
rect 3550 20417 3568 20451
rect 3516 20408 3568 20417
rect 5448 20476 5500 20528
rect 5080 20451 5132 20460
rect 5080 20417 5114 20451
rect 5114 20417 5132 20451
rect 5080 20408 5132 20417
rect 6736 20451 6788 20460
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 7104 20408 7156 20460
rect 8576 20476 8628 20528
rect 9588 20476 9640 20528
rect 11428 20544 11480 20596
rect 14740 20544 14792 20596
rect 15384 20544 15436 20596
rect 15660 20587 15712 20596
rect 15660 20553 15669 20587
rect 15669 20553 15703 20587
rect 15703 20553 15712 20587
rect 15660 20544 15712 20553
rect 15844 20544 15896 20596
rect 10324 20476 10376 20528
rect 12716 20476 12768 20528
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 9864 20408 9916 20460
rect 11244 20408 11296 20460
rect 11336 20408 11388 20460
rect 15200 20476 15252 20528
rect 16212 20476 16264 20528
rect 16488 20476 16540 20528
rect 14004 20408 14056 20460
rect 14464 20408 14516 20460
rect 14740 20408 14792 20460
rect 6460 20383 6512 20392
rect 6460 20349 6469 20383
rect 6469 20349 6503 20383
rect 6503 20349 6512 20383
rect 6460 20340 6512 20349
rect 15568 20383 15620 20392
rect 15568 20349 15577 20383
rect 15577 20349 15611 20383
rect 15611 20349 15620 20383
rect 15568 20340 15620 20349
rect 16028 20340 16080 20392
rect 16764 20408 16816 20460
rect 17224 20340 17276 20392
rect 19984 20544 20036 20596
rect 18972 20451 19024 20460
rect 18972 20417 18990 20451
rect 18990 20417 19024 20451
rect 18972 20408 19024 20417
rect 19800 20451 19852 20460
rect 19800 20417 19809 20451
rect 19809 20417 19843 20451
rect 19843 20417 19852 20451
rect 19800 20408 19852 20417
rect 20352 20544 20404 20596
rect 21272 20544 21324 20596
rect 20720 20476 20772 20528
rect 19248 20340 19300 20392
rect 19340 20383 19392 20392
rect 19340 20349 19349 20383
rect 19349 20349 19383 20383
rect 19383 20349 19392 20383
rect 19340 20340 19392 20349
rect 16948 20272 17000 20324
rect 4160 20204 4212 20256
rect 11520 20247 11572 20256
rect 11520 20213 11529 20247
rect 11529 20213 11563 20247
rect 11563 20213 11572 20247
rect 11520 20204 11572 20213
rect 15936 20204 15988 20256
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 22192 20204 22244 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 1350 20102 1402 20154
rect 1414 20102 1466 20154
rect 1478 20102 1530 20154
rect 1542 20102 1594 20154
rect 1606 20102 1658 20154
rect 4350 20102 4402 20154
rect 4414 20102 4466 20154
rect 4478 20102 4530 20154
rect 4542 20102 4594 20154
rect 4606 20102 4658 20154
rect 7350 20102 7402 20154
rect 7414 20102 7466 20154
rect 7478 20102 7530 20154
rect 7542 20102 7594 20154
rect 7606 20102 7658 20154
rect 10350 20102 10402 20154
rect 10414 20102 10466 20154
rect 10478 20102 10530 20154
rect 10542 20102 10594 20154
rect 10606 20102 10658 20154
rect 13350 20102 13402 20154
rect 13414 20102 13466 20154
rect 13478 20102 13530 20154
rect 13542 20102 13594 20154
rect 13606 20102 13658 20154
rect 16350 20102 16402 20154
rect 16414 20102 16466 20154
rect 16478 20102 16530 20154
rect 16542 20102 16594 20154
rect 16606 20102 16658 20154
rect 19350 20102 19402 20154
rect 19414 20102 19466 20154
rect 19478 20102 19530 20154
rect 19542 20102 19594 20154
rect 19606 20102 19658 20154
rect 22350 20102 22402 20154
rect 22414 20102 22466 20154
rect 22478 20102 22530 20154
rect 22542 20102 22594 20154
rect 22606 20102 22658 20154
rect 7196 20000 7248 20052
rect 8760 20000 8812 20052
rect 9680 20000 9732 20052
rect 11704 20000 11756 20052
rect 13912 20000 13964 20052
rect 16120 20043 16172 20052
rect 16120 20009 16129 20043
rect 16129 20009 16163 20043
rect 16163 20009 16172 20043
rect 16120 20000 16172 20009
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 18880 20000 18932 20052
rect 19248 20000 19300 20052
rect 19708 20000 19760 20052
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 9496 19864 9548 19873
rect 11520 19932 11572 19984
rect 10784 19907 10836 19916
rect 10784 19873 10793 19907
rect 10793 19873 10827 19907
rect 10827 19873 10836 19907
rect 10784 19864 10836 19873
rect 11152 19864 11204 19916
rect 6644 19796 6696 19848
rect 9404 19796 9456 19848
rect 11244 19796 11296 19848
rect 14372 19864 14424 19916
rect 15384 19864 15436 19916
rect 17500 19864 17552 19916
rect 17684 19864 17736 19916
rect 18972 19864 19024 19916
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16212 19796 16264 19848
rect 18604 19796 18656 19848
rect 19156 19796 19208 19848
rect 22836 19839 22888 19848
rect 22836 19805 22845 19839
rect 22845 19805 22879 19839
rect 22879 19805 22888 19839
rect 22836 19796 22888 19805
rect 22744 19728 22796 19780
rect 23020 19796 23072 19848
rect 23756 19796 23808 19848
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 21824 19660 21876 19712
rect 23112 19703 23164 19712
rect 23112 19669 23121 19703
rect 23121 19669 23155 19703
rect 23155 19669 23164 19703
rect 23112 19660 23164 19669
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 23664 19660 23716 19712
rect 2850 19558 2902 19610
rect 2914 19558 2966 19610
rect 2978 19558 3030 19610
rect 3042 19558 3094 19610
rect 3106 19558 3158 19610
rect 5850 19558 5902 19610
rect 5914 19558 5966 19610
rect 5978 19558 6030 19610
rect 6042 19558 6094 19610
rect 6106 19558 6158 19610
rect 8850 19558 8902 19610
rect 8914 19558 8966 19610
rect 8978 19558 9030 19610
rect 9042 19558 9094 19610
rect 9106 19558 9158 19610
rect 11850 19558 11902 19610
rect 11914 19558 11966 19610
rect 11978 19558 12030 19610
rect 12042 19558 12094 19610
rect 12106 19558 12158 19610
rect 14850 19558 14902 19610
rect 14914 19558 14966 19610
rect 14978 19558 15030 19610
rect 15042 19558 15094 19610
rect 15106 19558 15158 19610
rect 17850 19558 17902 19610
rect 17914 19558 17966 19610
rect 17978 19558 18030 19610
rect 18042 19558 18094 19610
rect 18106 19558 18158 19610
rect 20850 19558 20902 19610
rect 20914 19558 20966 19610
rect 20978 19558 21030 19610
rect 21042 19558 21094 19610
rect 21106 19558 21158 19610
rect 23850 19558 23902 19610
rect 23914 19558 23966 19610
rect 23978 19558 24030 19610
rect 24042 19558 24094 19610
rect 24106 19558 24158 19610
rect 9404 19499 9456 19508
rect 9404 19465 9413 19499
rect 9413 19465 9447 19499
rect 9447 19465 9456 19499
rect 9404 19456 9456 19465
rect 11612 19456 11664 19508
rect 13268 19456 13320 19508
rect 15292 19456 15344 19508
rect 16948 19456 17000 19508
rect 5632 19388 5684 19440
rect 3516 19363 3568 19372
rect 3516 19329 3550 19363
rect 3550 19329 3568 19363
rect 3516 19320 3568 19329
rect 1216 19116 1268 19168
rect 5264 19295 5316 19304
rect 5264 19261 5273 19295
rect 5273 19261 5307 19295
rect 5307 19261 5316 19295
rect 5264 19252 5316 19261
rect 6644 19320 6696 19372
rect 7012 19320 7064 19372
rect 23112 19388 23164 19440
rect 9680 19320 9732 19372
rect 11060 19320 11112 19372
rect 13912 19320 13964 19372
rect 16212 19320 16264 19372
rect 17684 19320 17736 19372
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 20720 19363 20772 19372
rect 20720 19329 20729 19363
rect 20729 19329 20763 19363
rect 20763 19329 20772 19363
rect 20720 19320 20772 19329
rect 21272 19320 21324 19372
rect 6092 19252 6144 19304
rect 6552 19252 6604 19304
rect 7104 19252 7156 19304
rect 9312 19252 9364 19304
rect 10692 19252 10744 19304
rect 10876 19252 10928 19304
rect 6460 19184 6512 19236
rect 10232 19184 10284 19236
rect 12348 19184 12400 19236
rect 14188 19252 14240 19304
rect 18788 19252 18840 19304
rect 19800 19252 19852 19304
rect 22928 19252 22980 19304
rect 23112 19295 23164 19304
rect 23112 19261 23121 19295
rect 23121 19261 23155 19295
rect 23155 19261 23164 19295
rect 23112 19252 23164 19261
rect 13728 19184 13780 19236
rect 15660 19184 15712 19236
rect 19892 19184 19944 19236
rect 23480 19184 23532 19236
rect 4160 19116 4212 19168
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 5448 19159 5500 19168
rect 5448 19125 5457 19159
rect 5457 19125 5491 19159
rect 5491 19125 5500 19159
rect 5448 19116 5500 19125
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 12716 19116 12768 19168
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 19708 19116 19760 19168
rect 20444 19116 20496 19168
rect 22100 19116 22152 19168
rect 23572 19159 23624 19168
rect 23572 19125 23581 19159
rect 23581 19125 23615 19159
rect 23615 19125 23624 19159
rect 23572 19116 23624 19125
rect 1350 19014 1402 19066
rect 1414 19014 1466 19066
rect 1478 19014 1530 19066
rect 1542 19014 1594 19066
rect 1606 19014 1658 19066
rect 4350 19014 4402 19066
rect 4414 19014 4466 19066
rect 4478 19014 4530 19066
rect 4542 19014 4594 19066
rect 4606 19014 4658 19066
rect 7350 19014 7402 19066
rect 7414 19014 7466 19066
rect 7478 19014 7530 19066
rect 7542 19014 7594 19066
rect 7606 19014 7658 19066
rect 10350 19014 10402 19066
rect 10414 19014 10466 19066
rect 10478 19014 10530 19066
rect 10542 19014 10594 19066
rect 10606 19014 10658 19066
rect 13350 19014 13402 19066
rect 13414 19014 13466 19066
rect 13478 19014 13530 19066
rect 13542 19014 13594 19066
rect 13606 19014 13658 19066
rect 16350 19014 16402 19066
rect 16414 19014 16466 19066
rect 16478 19014 16530 19066
rect 16542 19014 16594 19066
rect 16606 19014 16658 19066
rect 19350 19014 19402 19066
rect 19414 19014 19466 19066
rect 19478 19014 19530 19066
rect 19542 19014 19594 19066
rect 19606 19014 19658 19066
rect 22350 19014 22402 19066
rect 22414 19014 22466 19066
rect 22478 19014 22530 19066
rect 22542 19014 22594 19066
rect 22606 19014 22658 19066
rect 3516 18912 3568 18964
rect 5632 18912 5684 18964
rect 7104 18955 7156 18964
rect 7104 18921 7113 18955
rect 7113 18921 7147 18955
rect 7147 18921 7156 18955
rect 7104 18912 7156 18921
rect 16120 18912 16172 18964
rect 388 18708 440 18760
rect 3608 18751 3660 18760
rect 3608 18717 3617 18751
rect 3617 18717 3651 18751
rect 3651 18717 3660 18751
rect 3608 18708 3660 18717
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 5080 18708 5132 18760
rect 4712 18640 4764 18692
rect 5264 18776 5316 18828
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 6276 18776 6328 18828
rect 6736 18776 6788 18828
rect 9680 18776 9732 18828
rect 10232 18776 10284 18828
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 6920 18708 6972 18760
rect 9496 18708 9548 18760
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 11704 18708 11756 18760
rect 13820 18776 13872 18828
rect 15292 18776 15344 18828
rect 13268 18708 13320 18760
rect 7748 18640 7800 18692
rect 8668 18640 8720 18692
rect 10692 18640 10744 18692
rect 10968 18640 11020 18692
rect 14464 18708 14516 18760
rect 15384 18708 15436 18760
rect 17408 18708 17460 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 19708 18819 19760 18828
rect 19708 18785 19717 18819
rect 19717 18785 19751 18819
rect 19751 18785 19760 18819
rect 19708 18776 19760 18785
rect 21364 18912 21416 18964
rect 22836 18912 22888 18964
rect 22928 18844 22980 18896
rect 20168 18819 20220 18828
rect 20168 18785 20177 18819
rect 20177 18785 20211 18819
rect 20211 18785 20220 18819
rect 20168 18776 20220 18785
rect 19340 18708 19392 18760
rect 19892 18708 19944 18760
rect 20444 18751 20496 18760
rect 20444 18717 20478 18751
rect 20478 18717 20496 18751
rect 20444 18708 20496 18717
rect 22100 18819 22152 18828
rect 22100 18785 22109 18819
rect 22109 18785 22143 18819
rect 22143 18785 22152 18819
rect 22100 18776 22152 18785
rect 22376 18776 22428 18828
rect 22744 18708 22796 18760
rect 16856 18640 16908 18692
rect 8760 18572 8812 18624
rect 9312 18572 9364 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 14648 18572 14700 18624
rect 14740 18572 14792 18624
rect 16028 18572 16080 18624
rect 18788 18640 18840 18692
rect 19984 18640 20036 18692
rect 18236 18572 18288 18624
rect 20260 18572 20312 18624
rect 22100 18572 22152 18624
rect 22284 18572 22336 18624
rect 22744 18572 22796 18624
rect 24308 18572 24360 18624
rect 2850 18470 2902 18522
rect 2914 18470 2966 18522
rect 2978 18470 3030 18522
rect 3042 18470 3094 18522
rect 3106 18470 3158 18522
rect 5850 18470 5902 18522
rect 5914 18470 5966 18522
rect 5978 18470 6030 18522
rect 6042 18470 6094 18522
rect 6106 18470 6158 18522
rect 8850 18470 8902 18522
rect 8914 18470 8966 18522
rect 8978 18470 9030 18522
rect 9042 18470 9094 18522
rect 9106 18470 9158 18522
rect 11850 18470 11902 18522
rect 11914 18470 11966 18522
rect 11978 18470 12030 18522
rect 12042 18470 12094 18522
rect 12106 18470 12158 18522
rect 14850 18470 14902 18522
rect 14914 18470 14966 18522
rect 14978 18470 15030 18522
rect 15042 18470 15094 18522
rect 15106 18470 15158 18522
rect 17850 18470 17902 18522
rect 17914 18470 17966 18522
rect 17978 18470 18030 18522
rect 18042 18470 18094 18522
rect 18106 18470 18158 18522
rect 20850 18470 20902 18522
rect 20914 18470 20966 18522
rect 20978 18470 21030 18522
rect 21042 18470 21094 18522
rect 21106 18470 21158 18522
rect 23850 18470 23902 18522
rect 23914 18470 23966 18522
rect 23978 18470 24030 18522
rect 24042 18470 24094 18522
rect 24106 18470 24158 18522
rect 3608 18368 3660 18420
rect 5448 18368 5500 18420
rect 7196 18368 7248 18420
rect 8760 18411 8812 18420
rect 8760 18377 8769 18411
rect 8769 18377 8803 18411
rect 8803 18377 8812 18411
rect 8760 18368 8812 18377
rect 3792 18300 3844 18352
rect 5080 18343 5132 18352
rect 5080 18309 5089 18343
rect 5089 18309 5123 18343
rect 5123 18309 5132 18343
rect 5080 18300 5132 18309
rect 6644 18300 6696 18352
rect 7012 18300 7064 18352
rect 8668 18300 8720 18352
rect 10876 18368 10928 18420
rect 10232 18300 10284 18352
rect 14464 18368 14516 18420
rect 14648 18368 14700 18420
rect 12532 18300 12584 18352
rect 15384 18368 15436 18420
rect 16028 18411 16080 18420
rect 16028 18377 16037 18411
rect 16037 18377 16071 18411
rect 16071 18377 16080 18411
rect 16028 18368 16080 18377
rect 18512 18368 18564 18420
rect 6368 18232 6420 18284
rect 6460 18232 6512 18284
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 9312 18275 9364 18284
rect 9312 18241 9321 18275
rect 9321 18241 9355 18275
rect 9355 18241 9364 18275
rect 9312 18232 9364 18241
rect 9680 18232 9732 18284
rect 11152 18232 11204 18284
rect 12716 18232 12768 18284
rect 14464 18275 14516 18284
rect 14464 18241 14482 18275
rect 14482 18241 14516 18275
rect 14464 18232 14516 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 5172 18164 5224 18173
rect 5264 18096 5316 18148
rect 6920 18164 6972 18216
rect 11704 18164 11756 18216
rect 13912 18164 13964 18216
rect 15844 18232 15896 18284
rect 16672 18275 16724 18284
rect 16672 18241 16681 18275
rect 16681 18241 16715 18275
rect 16715 18241 16724 18275
rect 16672 18232 16724 18241
rect 18788 18275 18840 18284
rect 18788 18241 18797 18275
rect 18797 18241 18831 18275
rect 18831 18241 18840 18275
rect 18788 18232 18840 18241
rect 19708 18300 19760 18352
rect 19984 18411 20036 18420
rect 19984 18377 19993 18411
rect 19993 18377 20027 18411
rect 20027 18377 20036 18411
rect 19984 18368 20036 18377
rect 22652 18368 22704 18420
rect 4160 18028 4212 18080
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 7104 18028 7156 18080
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 11980 18071 12032 18080
rect 11980 18037 11989 18071
rect 11989 18037 12023 18071
rect 12023 18037 12032 18071
rect 11980 18028 12032 18037
rect 12440 18028 12492 18080
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15384 18164 15436 18216
rect 16120 18207 16172 18216
rect 16120 18173 16129 18207
rect 16129 18173 16163 18207
rect 16163 18173 16172 18207
rect 16120 18164 16172 18173
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 18512 18207 18564 18216
rect 14924 18096 14976 18148
rect 17316 18096 17368 18148
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 18696 18207 18748 18216
rect 18696 18173 18714 18207
rect 18714 18173 18748 18207
rect 18696 18164 18748 18173
rect 19156 18096 19208 18148
rect 20168 18232 20220 18284
rect 20352 18275 20404 18284
rect 20352 18241 20386 18275
rect 20386 18241 20404 18275
rect 20352 18232 20404 18241
rect 19892 18164 19944 18216
rect 22652 18275 22704 18284
rect 22652 18241 22670 18275
rect 22670 18241 22704 18275
rect 22652 18232 22704 18241
rect 22008 18096 22060 18148
rect 22928 18164 22980 18216
rect 23480 18207 23532 18216
rect 23480 18173 23489 18207
rect 23489 18173 23523 18207
rect 23523 18173 23532 18207
rect 23480 18164 23532 18173
rect 22560 18028 22612 18080
rect 22928 18028 22980 18080
rect 23112 18096 23164 18148
rect 1350 17926 1402 17978
rect 1414 17926 1466 17978
rect 1478 17926 1530 17978
rect 1542 17926 1594 17978
rect 1606 17926 1658 17978
rect 4350 17926 4402 17978
rect 4414 17926 4466 17978
rect 4478 17926 4530 17978
rect 4542 17926 4594 17978
rect 4606 17926 4658 17978
rect 7350 17926 7402 17978
rect 7414 17926 7466 17978
rect 7478 17926 7530 17978
rect 7542 17926 7594 17978
rect 7606 17926 7658 17978
rect 10350 17926 10402 17978
rect 10414 17926 10466 17978
rect 10478 17926 10530 17978
rect 10542 17926 10594 17978
rect 10606 17926 10658 17978
rect 13350 17926 13402 17978
rect 13414 17926 13466 17978
rect 13478 17926 13530 17978
rect 13542 17926 13594 17978
rect 13606 17926 13658 17978
rect 16350 17926 16402 17978
rect 16414 17926 16466 17978
rect 16478 17926 16530 17978
rect 16542 17926 16594 17978
rect 16606 17926 16658 17978
rect 19350 17926 19402 17978
rect 19414 17926 19466 17978
rect 19478 17926 19530 17978
rect 19542 17926 19594 17978
rect 19606 17926 19658 17978
rect 22350 17926 22402 17978
rect 22414 17926 22466 17978
rect 22478 17926 22530 17978
rect 22542 17926 22594 17978
rect 22606 17926 22658 17978
rect 6920 17824 6972 17876
rect 7748 17824 7800 17876
rect 11060 17824 11112 17876
rect 14188 17824 14240 17876
rect 14556 17824 14608 17876
rect 15292 17824 15344 17876
rect 17684 17824 17736 17876
rect 19708 17824 19760 17876
rect 23112 17867 23164 17876
rect 23112 17833 23121 17867
rect 23121 17833 23155 17867
rect 23155 17833 23164 17867
rect 23112 17824 23164 17833
rect 17500 17756 17552 17808
rect 9588 17688 9640 17740
rect 10232 17688 10284 17740
rect 10692 17688 10744 17740
rect 10876 17688 10928 17740
rect 11428 17688 11480 17740
rect 11704 17688 11756 17740
rect 4160 17620 4212 17672
rect 5632 17595 5684 17604
rect 5632 17561 5666 17595
rect 5666 17561 5684 17595
rect 5632 17552 5684 17561
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 7196 17620 7248 17672
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 9864 17620 9916 17672
rect 11336 17620 11388 17672
rect 11980 17620 12032 17672
rect 14096 17620 14148 17672
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 14648 17620 14700 17672
rect 17408 17620 17460 17672
rect 7748 17552 7800 17604
rect 8668 17484 8720 17536
rect 14832 17595 14884 17604
rect 14832 17561 14866 17595
rect 14866 17561 14884 17595
rect 14832 17552 14884 17561
rect 16948 17552 17000 17604
rect 11060 17527 11112 17536
rect 11060 17493 11069 17527
rect 11069 17493 11103 17527
rect 11103 17493 11112 17527
rect 11060 17484 11112 17493
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 13820 17484 13872 17536
rect 18236 17731 18288 17740
rect 18236 17697 18245 17731
rect 18245 17697 18279 17731
rect 18279 17697 18288 17731
rect 18236 17688 18288 17697
rect 17684 17620 17736 17672
rect 18512 17620 18564 17672
rect 19248 17688 19300 17740
rect 21640 17688 21692 17740
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 20628 17663 20680 17672
rect 20628 17629 20637 17663
rect 20637 17629 20671 17663
rect 20671 17629 20680 17663
rect 20628 17620 20680 17629
rect 18696 17552 18748 17604
rect 20168 17552 20220 17604
rect 20260 17552 20312 17604
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 20536 17484 20588 17536
rect 21824 17552 21876 17604
rect 22284 17620 22336 17672
rect 22744 17552 22796 17604
rect 22100 17484 22152 17536
rect 23388 17484 23440 17536
rect 2850 17382 2902 17434
rect 2914 17382 2966 17434
rect 2978 17382 3030 17434
rect 3042 17382 3094 17434
rect 3106 17382 3158 17434
rect 5850 17382 5902 17434
rect 5914 17382 5966 17434
rect 5978 17382 6030 17434
rect 6042 17382 6094 17434
rect 6106 17382 6158 17434
rect 8850 17382 8902 17434
rect 8914 17382 8966 17434
rect 8978 17382 9030 17434
rect 9042 17382 9094 17434
rect 9106 17382 9158 17434
rect 11850 17382 11902 17434
rect 11914 17382 11966 17434
rect 11978 17382 12030 17434
rect 12042 17382 12094 17434
rect 12106 17382 12158 17434
rect 14850 17382 14902 17434
rect 14914 17382 14966 17434
rect 14978 17382 15030 17434
rect 15042 17382 15094 17434
rect 15106 17382 15158 17434
rect 17850 17382 17902 17434
rect 17914 17382 17966 17434
rect 17978 17382 18030 17434
rect 18042 17382 18094 17434
rect 18106 17382 18158 17434
rect 20850 17382 20902 17434
rect 20914 17382 20966 17434
rect 20978 17382 21030 17434
rect 21042 17382 21094 17434
rect 21106 17382 21158 17434
rect 23850 17382 23902 17434
rect 23914 17382 23966 17434
rect 23978 17382 24030 17434
rect 24042 17382 24094 17434
rect 24106 17382 24158 17434
rect 5264 17280 5316 17332
rect 5724 17280 5776 17332
rect 6828 17280 6880 17332
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 6552 17212 6604 17264
rect 10784 17280 10836 17332
rect 11336 17323 11388 17332
rect 11336 17289 11345 17323
rect 11345 17289 11379 17323
rect 11379 17289 11388 17323
rect 11336 17280 11388 17289
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 15384 17280 15436 17332
rect 16856 17280 16908 17332
rect 9680 17212 9732 17264
rect 5540 17144 5592 17196
rect 5632 17144 5684 17196
rect 4252 17008 4304 17060
rect 5724 17008 5776 17060
rect 6460 17076 6512 17128
rect 8392 17076 8444 17128
rect 6552 17008 6604 17060
rect 6736 17008 6788 17060
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 5448 16940 5500 16992
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 10232 17187 10284 17196
rect 10232 17153 10266 17187
rect 10266 17153 10284 17187
rect 10232 17144 10284 17153
rect 11704 17212 11756 17264
rect 12348 17212 12400 17264
rect 13544 17255 13596 17264
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 12716 17144 12768 17196
rect 13544 17221 13578 17255
rect 13578 17221 13596 17255
rect 13544 17212 13596 17221
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 17776 17280 17828 17332
rect 19892 17280 19944 17332
rect 20352 17280 20404 17332
rect 22284 17280 22336 17332
rect 23480 17280 23532 17332
rect 17408 17212 17460 17264
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 18604 17212 18656 17264
rect 20628 17212 20680 17264
rect 20536 17144 20588 17196
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 21272 17144 21324 17196
rect 23204 17212 23256 17264
rect 9496 17076 9548 17128
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 9864 17076 9916 17128
rect 14556 17008 14608 17060
rect 15660 17051 15712 17060
rect 15660 17017 15669 17051
rect 15669 17017 15703 17051
rect 15703 17017 15712 17051
rect 15660 17008 15712 17017
rect 19064 17008 19116 17060
rect 10140 16940 10192 16992
rect 1350 16838 1402 16890
rect 1414 16838 1466 16890
rect 1478 16838 1530 16890
rect 1542 16838 1594 16890
rect 1606 16838 1658 16890
rect 4350 16838 4402 16890
rect 4414 16838 4466 16890
rect 4478 16838 4530 16890
rect 4542 16838 4594 16890
rect 4606 16838 4658 16890
rect 7350 16838 7402 16890
rect 7414 16838 7466 16890
rect 7478 16838 7530 16890
rect 7542 16838 7594 16890
rect 7606 16838 7658 16890
rect 10350 16838 10402 16890
rect 10414 16838 10466 16890
rect 10478 16838 10530 16890
rect 10542 16838 10594 16890
rect 10606 16838 10658 16890
rect 13350 16838 13402 16890
rect 13414 16838 13466 16890
rect 13478 16838 13530 16890
rect 13542 16838 13594 16890
rect 13606 16838 13658 16890
rect 16350 16838 16402 16890
rect 16414 16838 16466 16890
rect 16478 16838 16530 16890
rect 16542 16838 16594 16890
rect 16606 16838 16658 16890
rect 19350 16838 19402 16890
rect 19414 16838 19466 16890
rect 19478 16838 19530 16890
rect 19542 16838 19594 16890
rect 19606 16838 19658 16890
rect 22350 16838 22402 16890
rect 22414 16838 22466 16890
rect 22478 16838 22530 16890
rect 22542 16838 22594 16890
rect 22606 16838 22658 16890
rect 6644 16668 6696 16720
rect 3884 16600 3936 16652
rect 5724 16600 5776 16652
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 1308 16396 1360 16448
rect 2780 16532 2832 16584
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 6828 16736 6880 16788
rect 9772 16736 9824 16788
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 11428 16736 11480 16788
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 18788 16736 18840 16788
rect 20444 16736 20496 16788
rect 22100 16736 22152 16788
rect 9496 16668 9548 16720
rect 7196 16600 7248 16652
rect 8024 16532 8076 16584
rect 9588 16532 9640 16584
rect 9680 16532 9732 16584
rect 11060 16600 11112 16652
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 2504 16507 2556 16516
rect 2504 16473 2538 16507
rect 2538 16473 2556 16507
rect 2504 16464 2556 16473
rect 4252 16396 4304 16448
rect 4436 16396 4488 16448
rect 12716 16464 12768 16516
rect 14372 16532 14424 16584
rect 16856 16532 16908 16584
rect 17684 16532 17736 16584
rect 19064 16600 19116 16652
rect 21180 16600 21232 16652
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 21088 16575 21140 16584
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 14464 16507 14516 16516
rect 14464 16473 14473 16507
rect 14473 16473 14507 16507
rect 14507 16473 14516 16507
rect 14464 16464 14516 16473
rect 18512 16464 18564 16516
rect 15936 16396 15988 16448
rect 21732 16600 21784 16652
rect 22192 16643 22244 16652
rect 22192 16609 22201 16643
rect 22201 16609 22235 16643
rect 22235 16609 22244 16643
rect 22192 16600 22244 16609
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 23480 16643 23532 16652
rect 23480 16609 23489 16643
rect 23489 16609 23523 16643
rect 23523 16609 23532 16643
rect 23480 16600 23532 16609
rect 23020 16396 23072 16448
rect 2850 16294 2902 16346
rect 2914 16294 2966 16346
rect 2978 16294 3030 16346
rect 3042 16294 3094 16346
rect 3106 16294 3158 16346
rect 5850 16294 5902 16346
rect 5914 16294 5966 16346
rect 5978 16294 6030 16346
rect 6042 16294 6094 16346
rect 6106 16294 6158 16346
rect 8850 16294 8902 16346
rect 8914 16294 8966 16346
rect 8978 16294 9030 16346
rect 9042 16294 9094 16346
rect 9106 16294 9158 16346
rect 11850 16294 11902 16346
rect 11914 16294 11966 16346
rect 11978 16294 12030 16346
rect 12042 16294 12094 16346
rect 12106 16294 12158 16346
rect 14850 16294 14902 16346
rect 14914 16294 14966 16346
rect 14978 16294 15030 16346
rect 15042 16294 15094 16346
rect 15106 16294 15158 16346
rect 17850 16294 17902 16346
rect 17914 16294 17966 16346
rect 17978 16294 18030 16346
rect 18042 16294 18094 16346
rect 18106 16294 18158 16346
rect 20850 16294 20902 16346
rect 20914 16294 20966 16346
rect 20978 16294 21030 16346
rect 21042 16294 21094 16346
rect 21106 16294 21158 16346
rect 23850 16294 23902 16346
rect 23914 16294 23966 16346
rect 23978 16294 24030 16346
rect 24042 16294 24094 16346
rect 24106 16294 24158 16346
rect 2504 16192 2556 16244
rect 2780 16192 2832 16244
rect 3884 16235 3936 16244
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 3884 16192 3936 16201
rect 4436 16235 4488 16244
rect 4436 16201 4445 16235
rect 4445 16201 4479 16235
rect 4479 16201 4488 16235
rect 4436 16192 4488 16201
rect 6460 16192 6512 16244
rect 15936 16235 15988 16244
rect 15936 16201 15945 16235
rect 15945 16201 15979 16235
rect 15979 16201 15988 16235
rect 15936 16192 15988 16201
rect 20628 16192 20680 16244
rect 756 16056 808 16108
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2872 16124 2924 16176
rect 5264 16124 5316 16176
rect 6276 16124 6328 16176
rect 3516 15920 3568 15972
rect 4160 15852 4212 15904
rect 5632 16056 5684 16108
rect 16028 16124 16080 16176
rect 18788 16124 18840 16176
rect 20720 16124 20772 16176
rect 22192 16124 22244 16176
rect 8300 16056 8352 16108
rect 11888 16056 11940 16108
rect 14004 16056 14056 16108
rect 15568 16056 15620 16108
rect 16304 16056 16356 16108
rect 4712 15988 4764 16040
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 6644 15988 6696 16040
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 12992 15988 13044 16040
rect 16212 15988 16264 16040
rect 9956 15920 10008 15972
rect 13268 15920 13320 15972
rect 16764 15920 16816 15972
rect 17684 15920 17736 15972
rect 18604 16031 18656 16040
rect 18604 15997 18613 16031
rect 18613 15997 18647 16031
rect 18647 15997 18656 16031
rect 18604 15988 18656 15997
rect 21088 16056 21140 16108
rect 5540 15852 5592 15904
rect 7932 15852 7984 15904
rect 10968 15852 11020 15904
rect 11704 15852 11756 15904
rect 12808 15852 12860 15904
rect 15108 15852 15160 15904
rect 15384 15852 15436 15904
rect 18972 15852 19024 15904
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 20720 15988 20772 16040
rect 21916 15988 21968 16040
rect 21180 15920 21232 15972
rect 21364 15920 21416 15972
rect 21824 15920 21876 15972
rect 20628 15852 20680 15904
rect 20812 15852 20864 15904
rect 23664 15852 23716 15904
rect 1350 15750 1402 15802
rect 1414 15750 1466 15802
rect 1478 15750 1530 15802
rect 1542 15750 1594 15802
rect 1606 15750 1658 15802
rect 4350 15750 4402 15802
rect 4414 15750 4466 15802
rect 4478 15750 4530 15802
rect 4542 15750 4594 15802
rect 4606 15750 4658 15802
rect 7350 15750 7402 15802
rect 7414 15750 7466 15802
rect 7478 15750 7530 15802
rect 7542 15750 7594 15802
rect 7606 15750 7658 15802
rect 10350 15750 10402 15802
rect 10414 15750 10466 15802
rect 10478 15750 10530 15802
rect 10542 15750 10594 15802
rect 10606 15750 10658 15802
rect 13350 15750 13402 15802
rect 13414 15750 13466 15802
rect 13478 15750 13530 15802
rect 13542 15750 13594 15802
rect 13606 15750 13658 15802
rect 16350 15750 16402 15802
rect 16414 15750 16466 15802
rect 16478 15750 16530 15802
rect 16542 15750 16594 15802
rect 16606 15750 16658 15802
rect 19350 15750 19402 15802
rect 19414 15750 19466 15802
rect 19478 15750 19530 15802
rect 19542 15750 19594 15802
rect 19606 15750 19658 15802
rect 22350 15750 22402 15802
rect 22414 15750 22466 15802
rect 22478 15750 22530 15802
rect 22542 15750 22594 15802
rect 22606 15750 22658 15802
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 2228 15580 2280 15632
rect 6276 15648 6328 15700
rect 9680 15648 9732 15700
rect 7932 15580 7984 15632
rect 8116 15580 8168 15632
rect 10140 15580 10192 15632
rect 2780 15512 2832 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 3516 15444 3568 15496
rect 4160 15512 4212 15564
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 8300 15512 8352 15564
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 14096 15648 14148 15700
rect 11520 15580 11572 15632
rect 17500 15648 17552 15700
rect 11428 15512 11480 15564
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 12348 15555 12400 15564
rect 12348 15521 12357 15555
rect 12357 15521 12391 15555
rect 12391 15521 12400 15555
rect 12348 15512 12400 15521
rect 16672 15512 16724 15564
rect 17776 15623 17828 15632
rect 17776 15589 17785 15623
rect 17785 15589 17819 15623
rect 17819 15589 17828 15623
rect 17776 15580 17828 15589
rect 19248 15580 19300 15632
rect 20720 15691 20772 15700
rect 20720 15657 20729 15691
rect 20729 15657 20763 15691
rect 20763 15657 20772 15691
rect 20720 15648 20772 15657
rect 21272 15648 21324 15700
rect 23296 15648 23348 15700
rect 22284 15623 22336 15632
rect 22284 15589 22293 15623
rect 22293 15589 22327 15623
rect 22327 15589 22336 15623
rect 22284 15580 22336 15589
rect 22836 15580 22888 15632
rect 17040 15512 17092 15564
rect 17215 15555 17267 15564
rect 17215 15521 17223 15555
rect 17223 15521 17257 15555
rect 17257 15521 17267 15555
rect 17215 15512 17267 15521
rect 17500 15555 17552 15564
rect 17500 15521 17509 15555
rect 17509 15521 17543 15555
rect 17543 15521 17552 15555
rect 17500 15512 17552 15521
rect 18604 15512 18656 15564
rect 22192 15512 22244 15564
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 5080 15487 5132 15496
rect 5080 15453 5114 15487
rect 5114 15453 5132 15487
rect 5080 15444 5132 15453
rect 7748 15444 7800 15496
rect 9680 15444 9732 15496
rect 9956 15487 10008 15496
rect 9956 15453 9965 15487
rect 9965 15453 9999 15487
rect 9999 15453 10008 15487
rect 9956 15444 10008 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 14740 15444 14792 15496
rect 15108 15487 15160 15496
rect 15108 15453 15142 15487
rect 15142 15453 15160 15487
rect 15108 15444 15160 15453
rect 17408 15487 17460 15512
rect 17408 15460 17426 15487
rect 17426 15460 17460 15487
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 7012 15376 7064 15428
rect 7564 15376 7616 15428
rect 4160 15351 4212 15360
rect 4160 15317 4169 15351
rect 4169 15317 4203 15351
rect 4203 15317 4212 15351
rect 4160 15308 4212 15317
rect 4712 15308 4764 15360
rect 8116 15308 8168 15360
rect 8208 15351 8260 15360
rect 8208 15317 8217 15351
rect 8217 15317 8251 15351
rect 8251 15317 8260 15351
rect 8208 15308 8260 15317
rect 9588 15351 9640 15360
rect 9588 15317 9597 15351
rect 9597 15317 9631 15351
rect 9631 15317 9640 15351
rect 9588 15308 9640 15317
rect 10232 15308 10284 15360
rect 11336 15351 11388 15360
rect 11336 15317 11345 15351
rect 11345 15317 11379 15351
rect 11379 15317 11388 15351
rect 11336 15308 11388 15317
rect 12440 15376 12492 15428
rect 12900 15308 12952 15360
rect 13912 15308 13964 15360
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 19340 15487 19392 15496
rect 19340 15453 19349 15487
rect 19349 15453 19383 15487
rect 19383 15453 19392 15487
rect 19340 15444 19392 15453
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 21916 15487 21968 15496
rect 21916 15453 21934 15487
rect 21934 15453 21968 15487
rect 21916 15444 21968 15453
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 23020 15444 23072 15496
rect 23112 15487 23164 15496
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 19800 15376 19852 15428
rect 18788 15308 18840 15360
rect 21088 15376 21140 15428
rect 21456 15308 21508 15360
rect 2850 15206 2902 15258
rect 2914 15206 2966 15258
rect 2978 15206 3030 15258
rect 3042 15206 3094 15258
rect 3106 15206 3158 15258
rect 5850 15206 5902 15258
rect 5914 15206 5966 15258
rect 5978 15206 6030 15258
rect 6042 15206 6094 15258
rect 6106 15206 6158 15258
rect 8850 15206 8902 15258
rect 8914 15206 8966 15258
rect 8978 15206 9030 15258
rect 9042 15206 9094 15258
rect 9106 15206 9158 15258
rect 11850 15206 11902 15258
rect 11914 15206 11966 15258
rect 11978 15206 12030 15258
rect 12042 15206 12094 15258
rect 12106 15206 12158 15258
rect 14850 15206 14902 15258
rect 14914 15206 14966 15258
rect 14978 15206 15030 15258
rect 15042 15206 15094 15258
rect 15106 15206 15158 15258
rect 17850 15206 17902 15258
rect 17914 15206 17966 15258
rect 17978 15206 18030 15258
rect 18042 15206 18094 15258
rect 18106 15206 18158 15258
rect 20850 15206 20902 15258
rect 20914 15206 20966 15258
rect 20978 15206 21030 15258
rect 21042 15206 21094 15258
rect 21106 15206 21158 15258
rect 23850 15206 23902 15258
rect 23914 15206 23966 15258
rect 23978 15206 24030 15258
rect 24042 15206 24094 15258
rect 24106 15206 24158 15258
rect 4160 15104 4212 15156
rect 5264 15147 5316 15156
rect 5264 15113 5273 15147
rect 5273 15113 5307 15147
rect 5307 15113 5316 15147
rect 5264 15104 5316 15113
rect 4252 15036 4304 15088
rect 1216 14968 1268 15020
rect 2964 14968 3016 15020
rect 3332 14968 3384 15020
rect 4436 14968 4488 15020
rect 5448 15011 5500 15020
rect 5448 14977 5457 15011
rect 5457 14977 5491 15011
rect 5491 14977 5500 15011
rect 5448 14968 5500 14977
rect 7564 15104 7616 15156
rect 8208 15104 8260 15156
rect 9496 15104 9548 15156
rect 11244 15104 11296 15156
rect 12440 15104 12492 15156
rect 12900 15104 12952 15156
rect 13084 15104 13136 15156
rect 4252 14900 4304 14952
rect 4896 14900 4948 14952
rect 9404 14968 9456 15020
rect 11520 15036 11572 15088
rect 14004 15147 14056 15156
rect 14004 15113 14013 15147
rect 14013 15113 14047 15147
rect 14047 15113 14056 15147
rect 14004 15104 14056 15113
rect 6644 14832 6696 14884
rect 2688 14764 2740 14816
rect 2872 14764 2924 14816
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 8300 14832 8352 14884
rect 9128 14764 9180 14816
rect 10048 14968 10100 15020
rect 11336 14968 11388 15020
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 12716 15011 12768 15020
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 16120 15104 16172 15156
rect 16856 15104 16908 15156
rect 17408 15104 17460 15156
rect 18604 15104 18656 15156
rect 18788 15147 18840 15156
rect 18788 15113 18797 15147
rect 18797 15113 18831 15147
rect 18831 15113 18840 15147
rect 18788 15104 18840 15113
rect 18972 15104 19024 15156
rect 20444 15104 20496 15156
rect 21732 15104 21784 15156
rect 23388 15104 23440 15156
rect 14740 15036 14792 15088
rect 15108 15011 15160 15020
rect 15108 14977 15142 15011
rect 15142 14977 15160 15011
rect 15108 14968 15160 14977
rect 11244 14900 11296 14952
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13728 14943 13780 14952
rect 13728 14909 13737 14943
rect 13737 14909 13771 14943
rect 13771 14909 13780 14943
rect 13728 14900 13780 14909
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 16488 15036 16540 15088
rect 21824 15036 21876 15088
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 19984 14968 20036 15020
rect 20720 14968 20772 15020
rect 22928 15011 22980 15020
rect 22928 14977 22946 15011
rect 22946 14977 22980 15011
rect 22928 14968 22980 14977
rect 23296 14968 23348 15020
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 19340 14943 19392 14952
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 20996 14900 21048 14952
rect 21640 14900 21692 14952
rect 21916 14832 21968 14884
rect 11060 14764 11112 14816
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 14280 14764 14332 14816
rect 17224 14764 17276 14816
rect 20812 14807 20864 14816
rect 20812 14773 20821 14807
rect 20821 14773 20855 14807
rect 20855 14773 20864 14807
rect 20812 14764 20864 14773
rect 23020 14764 23072 14816
rect 1350 14662 1402 14714
rect 1414 14662 1466 14714
rect 1478 14662 1530 14714
rect 1542 14662 1594 14714
rect 1606 14662 1658 14714
rect 4350 14662 4402 14714
rect 4414 14662 4466 14714
rect 4478 14662 4530 14714
rect 4542 14662 4594 14714
rect 4606 14662 4658 14714
rect 7350 14662 7402 14714
rect 7414 14662 7466 14714
rect 7478 14662 7530 14714
rect 7542 14662 7594 14714
rect 7606 14662 7658 14714
rect 10350 14662 10402 14714
rect 10414 14662 10466 14714
rect 10478 14662 10530 14714
rect 10542 14662 10594 14714
rect 10606 14662 10658 14714
rect 13350 14662 13402 14714
rect 13414 14662 13466 14714
rect 13478 14662 13530 14714
rect 13542 14662 13594 14714
rect 13606 14662 13658 14714
rect 16350 14662 16402 14714
rect 16414 14662 16466 14714
rect 16478 14662 16530 14714
rect 16542 14662 16594 14714
rect 16606 14662 16658 14714
rect 19350 14662 19402 14714
rect 19414 14662 19466 14714
rect 19478 14662 19530 14714
rect 19542 14662 19594 14714
rect 19606 14662 19658 14714
rect 22350 14662 22402 14714
rect 22414 14662 22466 14714
rect 22478 14662 22530 14714
rect 22542 14662 22594 14714
rect 22606 14662 22658 14714
rect 2688 14424 2740 14476
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 2872 14356 2924 14408
rect 4896 14424 4948 14476
rect 4620 14356 4672 14408
rect 5724 14399 5776 14408
rect 5724 14365 5733 14399
rect 5733 14365 5767 14399
rect 5767 14365 5776 14399
rect 5724 14356 5776 14365
rect 6552 14356 6604 14408
rect 7380 14560 7432 14612
rect 7748 14560 7800 14612
rect 9404 14560 9456 14612
rect 10048 14560 10100 14612
rect 12900 14560 12952 14612
rect 13728 14560 13780 14612
rect 11796 14492 11848 14544
rect 12440 14492 12492 14544
rect 9128 14467 9180 14476
rect 9128 14433 9137 14467
rect 9137 14433 9171 14467
rect 9171 14433 9180 14467
rect 9128 14424 9180 14433
rect 9588 14424 9640 14476
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 7196 14356 7248 14408
rect 8760 14356 8812 14408
rect 14464 14560 14516 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 18236 14560 18288 14612
rect 14556 14492 14608 14544
rect 16948 14492 17000 14544
rect 756 14220 808 14272
rect 1860 14220 1912 14272
rect 9220 14288 9272 14340
rect 10232 14356 10284 14408
rect 14280 14424 14332 14476
rect 12808 14399 12860 14408
rect 12808 14365 12842 14399
rect 12842 14365 12860 14399
rect 12808 14356 12860 14365
rect 16028 14467 16080 14476
rect 16028 14433 16037 14467
rect 16037 14433 16071 14467
rect 16071 14433 16080 14467
rect 16028 14424 16080 14433
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 17040 14467 17092 14476
rect 17040 14433 17049 14467
rect 17049 14433 17083 14467
rect 17083 14433 17092 14467
rect 17040 14424 17092 14433
rect 18880 14560 18932 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 20996 14603 21048 14612
rect 20996 14569 21005 14603
rect 21005 14569 21039 14603
rect 21039 14569 21048 14603
rect 20996 14560 21048 14569
rect 23112 14560 23164 14612
rect 21916 14492 21968 14544
rect 3516 14220 3568 14272
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 6184 14220 6236 14272
rect 6920 14220 6972 14272
rect 7012 14220 7064 14272
rect 11520 14288 11572 14340
rect 11060 14220 11112 14272
rect 13820 14288 13872 14340
rect 14648 14288 14700 14340
rect 17224 14356 17276 14408
rect 20812 14356 20864 14408
rect 21824 14356 21876 14408
rect 22468 14356 22520 14408
rect 21456 14288 21508 14340
rect 15292 14220 15344 14272
rect 15844 14220 15896 14272
rect 23572 14263 23624 14272
rect 23572 14229 23581 14263
rect 23581 14229 23615 14263
rect 23615 14229 23624 14263
rect 23572 14220 23624 14229
rect 2850 14118 2902 14170
rect 2914 14118 2966 14170
rect 2978 14118 3030 14170
rect 3042 14118 3094 14170
rect 3106 14118 3158 14170
rect 5850 14118 5902 14170
rect 5914 14118 5966 14170
rect 5978 14118 6030 14170
rect 6042 14118 6094 14170
rect 6106 14118 6158 14170
rect 8850 14118 8902 14170
rect 8914 14118 8966 14170
rect 8978 14118 9030 14170
rect 9042 14118 9094 14170
rect 9106 14118 9158 14170
rect 11850 14118 11902 14170
rect 11914 14118 11966 14170
rect 11978 14118 12030 14170
rect 12042 14118 12094 14170
rect 12106 14118 12158 14170
rect 14850 14118 14902 14170
rect 14914 14118 14966 14170
rect 14978 14118 15030 14170
rect 15042 14118 15094 14170
rect 15106 14118 15158 14170
rect 17850 14118 17902 14170
rect 17914 14118 17966 14170
rect 17978 14118 18030 14170
rect 18042 14118 18094 14170
rect 18106 14118 18158 14170
rect 20850 14118 20902 14170
rect 20914 14118 20966 14170
rect 20978 14118 21030 14170
rect 21042 14118 21094 14170
rect 21106 14118 21158 14170
rect 23850 14118 23902 14170
rect 23914 14118 23966 14170
rect 23978 14118 24030 14170
rect 24042 14118 24094 14170
rect 24106 14118 24158 14170
rect 4068 14016 4120 14068
rect 4160 14016 4212 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 2780 13948 2832 14000
rect 3424 13948 3476 14000
rect 1676 13880 1728 13932
rect 1860 13923 1912 13932
rect 1860 13889 1894 13923
rect 1894 13889 1912 13923
rect 1860 13880 1912 13889
rect 3516 13923 3568 13932
rect 3516 13889 3550 13923
rect 3550 13889 3568 13923
rect 3516 13880 3568 13889
rect 4620 13787 4672 13796
rect 4620 13753 4629 13787
rect 4629 13753 4663 13787
rect 4663 13753 4672 13787
rect 4620 13744 4672 13753
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 8300 14016 8352 14068
rect 9220 14016 9272 14068
rect 9496 14016 9548 14068
rect 13728 14016 13780 14068
rect 15200 14059 15252 14068
rect 15200 14025 15209 14059
rect 15209 14025 15243 14059
rect 15243 14025 15252 14059
rect 15200 14016 15252 14025
rect 15844 14016 15896 14068
rect 22468 14016 22520 14068
rect 12532 13991 12584 14000
rect 12532 13957 12541 13991
rect 12541 13957 12575 13991
rect 12575 13957 12584 13991
rect 12532 13948 12584 13957
rect 15292 13948 15344 14000
rect 10692 13923 10744 13932
rect 10692 13889 10701 13923
rect 10701 13889 10735 13923
rect 10735 13889 10744 13923
rect 10692 13880 10744 13889
rect 13912 13880 13964 13932
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 20812 13948 20864 14000
rect 21088 13880 21140 13932
rect 22928 14016 22980 14068
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 5356 13812 5408 13864
rect 7932 13812 7984 13864
rect 4804 13744 4856 13796
rect 7840 13744 7892 13796
rect 4160 13676 4212 13728
rect 5264 13676 5316 13728
rect 6644 13676 6696 13728
rect 7104 13676 7156 13728
rect 8392 13855 8444 13864
rect 8392 13821 8426 13855
rect 8426 13821 8444 13855
rect 8392 13812 8444 13821
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 20720 13812 20772 13864
rect 21272 13812 21324 13864
rect 21916 13812 21968 13864
rect 17776 13744 17828 13796
rect 23020 13812 23072 13864
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 21364 13676 21416 13728
rect 22100 13676 22152 13728
rect 22836 13676 22888 13728
rect 1350 13574 1402 13626
rect 1414 13574 1466 13626
rect 1478 13574 1530 13626
rect 1542 13574 1594 13626
rect 1606 13574 1658 13626
rect 4350 13574 4402 13626
rect 4414 13574 4466 13626
rect 4478 13574 4530 13626
rect 4542 13574 4594 13626
rect 4606 13574 4658 13626
rect 7350 13574 7402 13626
rect 7414 13574 7466 13626
rect 7478 13574 7530 13626
rect 7542 13574 7594 13626
rect 7606 13574 7658 13626
rect 10350 13574 10402 13626
rect 10414 13574 10466 13626
rect 10478 13574 10530 13626
rect 10542 13574 10594 13626
rect 10606 13574 10658 13626
rect 13350 13574 13402 13626
rect 13414 13574 13466 13626
rect 13478 13574 13530 13626
rect 13542 13574 13594 13626
rect 13606 13574 13658 13626
rect 16350 13574 16402 13626
rect 16414 13574 16466 13626
rect 16478 13574 16530 13626
rect 16542 13574 16594 13626
rect 16606 13574 16658 13626
rect 19350 13574 19402 13626
rect 19414 13574 19466 13626
rect 19478 13574 19530 13626
rect 19542 13574 19594 13626
rect 19606 13574 19658 13626
rect 22350 13574 22402 13626
rect 22414 13574 22466 13626
rect 22478 13574 22530 13626
rect 22542 13574 22594 13626
rect 22606 13574 22658 13626
rect 1676 13472 1728 13524
rect 4252 13472 4304 13524
rect 4712 13472 4764 13524
rect 5724 13472 5776 13524
rect 7104 13472 7156 13524
rect 12440 13472 12492 13524
rect 13084 13472 13136 13524
rect 13268 13472 13320 13524
rect 20812 13515 20864 13524
rect 20812 13481 20821 13515
rect 20821 13481 20855 13515
rect 20855 13481 20864 13515
rect 20812 13472 20864 13481
rect 21088 13472 21140 13524
rect 23480 13472 23532 13524
rect 4160 13336 4212 13388
rect 4344 13336 4396 13388
rect 13176 13404 13228 13456
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 3884 13268 3936 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 1860 13200 1912 13252
rect 2596 13200 2648 13252
rect 3976 13132 4028 13184
rect 6184 13311 6236 13320
rect 6184 13277 6218 13311
rect 6218 13277 6236 13311
rect 6184 13268 6236 13277
rect 6644 13268 6696 13320
rect 8116 13336 8168 13388
rect 13728 13336 13780 13388
rect 7012 13268 7064 13320
rect 7840 13268 7892 13320
rect 8668 13268 8720 13320
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 12348 13311 12400 13320
rect 12348 13277 12357 13311
rect 12357 13277 12391 13311
rect 12391 13277 12400 13311
rect 12348 13268 12400 13277
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 14372 13268 14424 13320
rect 16212 13404 16264 13456
rect 16120 13336 16172 13388
rect 15936 13268 15988 13320
rect 18420 13336 18472 13388
rect 21640 13404 21692 13456
rect 20628 13336 20680 13388
rect 21364 13379 21416 13388
rect 21364 13345 21373 13379
rect 21373 13345 21407 13379
rect 21407 13345 21416 13379
rect 21364 13336 21416 13345
rect 8576 13200 8628 13252
rect 13176 13200 13228 13252
rect 15292 13200 15344 13252
rect 17500 13268 17552 13320
rect 20536 13268 20588 13320
rect 21548 13268 21600 13320
rect 21824 13268 21876 13320
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 18788 13200 18840 13252
rect 21180 13200 21232 13252
rect 21640 13200 21692 13252
rect 22192 13243 22244 13252
rect 22192 13209 22226 13243
rect 22226 13209 22244 13243
rect 22192 13200 22244 13209
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 11704 13132 11756 13184
rect 14740 13132 14792 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17132 13132 17184 13141
rect 17408 13175 17460 13184
rect 17408 13141 17417 13175
rect 17417 13141 17451 13175
rect 17451 13141 17460 13175
rect 17408 13132 17460 13141
rect 17592 13132 17644 13184
rect 19432 13132 19484 13184
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 20260 13175 20312 13184
rect 20260 13141 20269 13175
rect 20269 13141 20303 13175
rect 20303 13141 20312 13175
rect 20260 13132 20312 13141
rect 20628 13132 20680 13184
rect 21548 13132 21600 13184
rect 21916 13132 21968 13184
rect 22744 13132 22796 13184
rect 24308 13132 24360 13184
rect 2850 13030 2902 13082
rect 2914 13030 2966 13082
rect 2978 13030 3030 13082
rect 3042 13030 3094 13082
rect 3106 13030 3158 13082
rect 5850 13030 5902 13082
rect 5914 13030 5966 13082
rect 5978 13030 6030 13082
rect 6042 13030 6094 13082
rect 6106 13030 6158 13082
rect 8850 13030 8902 13082
rect 8914 13030 8966 13082
rect 8978 13030 9030 13082
rect 9042 13030 9094 13082
rect 9106 13030 9158 13082
rect 11850 13030 11902 13082
rect 11914 13030 11966 13082
rect 11978 13030 12030 13082
rect 12042 13030 12094 13082
rect 12106 13030 12158 13082
rect 14850 13030 14902 13082
rect 14914 13030 14966 13082
rect 14978 13030 15030 13082
rect 15042 13030 15094 13082
rect 15106 13030 15158 13082
rect 17850 13030 17902 13082
rect 17914 13030 17966 13082
rect 17978 13030 18030 13082
rect 18042 13030 18094 13082
rect 18106 13030 18158 13082
rect 20850 13030 20902 13082
rect 20914 13030 20966 13082
rect 20978 13030 21030 13082
rect 21042 13030 21094 13082
rect 21106 13030 21158 13082
rect 23850 13030 23902 13082
rect 23914 13030 23966 13082
rect 23978 13030 24030 13082
rect 24042 13030 24094 13082
rect 24106 13030 24158 13082
rect 1308 12928 1360 12980
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 3884 12928 3936 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 2688 12860 2740 12912
rect 2780 12860 2832 12912
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 4528 12792 4580 12844
rect 5540 12588 5592 12640
rect 7380 12928 7432 12980
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 8760 12860 8812 12912
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 8668 12656 8720 12708
rect 10140 12724 10192 12776
rect 11428 12928 11480 12980
rect 12348 12928 12400 12980
rect 12808 12928 12860 12980
rect 11336 12860 11388 12912
rect 11428 12792 11480 12844
rect 14740 12860 14792 12912
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 16028 12860 16080 12912
rect 17592 12835 17644 12844
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 17592 12792 17644 12801
rect 18788 12971 18840 12980
rect 18788 12937 18797 12971
rect 18797 12937 18831 12971
rect 18831 12937 18840 12971
rect 18788 12928 18840 12937
rect 19892 12928 19944 12980
rect 20536 12928 20588 12980
rect 20720 12928 20772 12980
rect 21180 12928 21232 12980
rect 23204 12928 23256 12980
rect 19156 12860 19208 12912
rect 21824 12860 21876 12912
rect 19432 12835 19484 12844
rect 19432 12801 19466 12835
rect 19466 12801 19484 12835
rect 19432 12792 19484 12801
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 22744 12835 22796 12844
rect 22744 12801 22753 12835
rect 22753 12801 22787 12835
rect 22787 12801 22796 12835
rect 22744 12792 22796 12801
rect 23296 12792 23348 12844
rect 11060 12724 11112 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 17776 12724 17828 12776
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 11796 12656 11848 12708
rect 18236 12656 18288 12708
rect 19156 12767 19208 12776
rect 19156 12733 19165 12767
rect 19165 12733 19199 12767
rect 19199 12733 19208 12767
rect 19156 12724 19208 12733
rect 20260 12724 20312 12776
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 21180 12656 21232 12708
rect 6644 12588 6696 12640
rect 9404 12588 9456 12640
rect 11520 12588 11572 12640
rect 12992 12588 13044 12640
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 19800 12588 19852 12640
rect 21364 12588 21416 12640
rect 22928 12724 22980 12776
rect 23480 12767 23532 12776
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 21916 12588 21968 12640
rect 22100 12588 22152 12640
rect 1350 12486 1402 12538
rect 1414 12486 1466 12538
rect 1478 12486 1530 12538
rect 1542 12486 1594 12538
rect 1606 12486 1658 12538
rect 4350 12486 4402 12538
rect 4414 12486 4466 12538
rect 4478 12486 4530 12538
rect 4542 12486 4594 12538
rect 4606 12486 4658 12538
rect 7350 12486 7402 12538
rect 7414 12486 7466 12538
rect 7478 12486 7530 12538
rect 7542 12486 7594 12538
rect 7606 12486 7658 12538
rect 10350 12486 10402 12538
rect 10414 12486 10466 12538
rect 10478 12486 10530 12538
rect 10542 12486 10594 12538
rect 10606 12486 10658 12538
rect 13350 12486 13402 12538
rect 13414 12486 13466 12538
rect 13478 12486 13530 12538
rect 13542 12486 13594 12538
rect 13606 12486 13658 12538
rect 16350 12486 16402 12538
rect 16414 12486 16466 12538
rect 16478 12486 16530 12538
rect 16542 12486 16594 12538
rect 16606 12486 16658 12538
rect 19350 12486 19402 12538
rect 19414 12486 19466 12538
rect 19478 12486 19530 12538
rect 19542 12486 19594 12538
rect 19606 12486 19658 12538
rect 22350 12486 22402 12538
rect 22414 12486 22466 12538
rect 22478 12486 22530 12538
rect 22542 12486 22594 12538
rect 22606 12486 22658 12538
rect 4252 12384 4304 12436
rect 10140 12384 10192 12436
rect 11428 12384 11480 12436
rect 11520 12384 11572 12436
rect 11796 12359 11848 12368
rect 11796 12325 11805 12359
rect 11805 12325 11839 12359
rect 11839 12325 11848 12359
rect 11796 12316 11848 12325
rect 11060 12248 11112 12300
rect 12348 12248 12400 12300
rect 388 12180 440 12232
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 8668 12180 8720 12232
rect 8760 12180 8812 12232
rect 9220 12180 9272 12232
rect 9404 12223 9456 12232
rect 9404 12189 9438 12223
rect 9438 12189 9456 12223
rect 9404 12180 9456 12189
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 11428 12223 11480 12232
rect 11428 12189 11446 12223
rect 11446 12189 11480 12223
rect 11428 12180 11480 12189
rect 12900 12180 12952 12232
rect 16028 12427 16080 12436
rect 16028 12393 16037 12427
rect 16037 12393 16071 12427
rect 16071 12393 16080 12427
rect 16028 12384 16080 12393
rect 16580 12384 16632 12436
rect 17776 12384 17828 12436
rect 18420 12384 18472 12436
rect 20720 12427 20772 12436
rect 20720 12393 20729 12427
rect 20729 12393 20763 12427
rect 20763 12393 20772 12427
rect 20720 12384 20772 12393
rect 22192 12384 22244 12436
rect 23296 12384 23348 12436
rect 16212 12248 16264 12300
rect 14096 12180 14148 12232
rect 14464 12180 14516 12232
rect 16856 12223 16908 12232
rect 16856 12189 16865 12223
rect 16865 12189 16899 12223
rect 16899 12189 16908 12223
rect 16856 12180 16908 12189
rect 17132 12223 17184 12232
rect 17132 12189 17166 12223
rect 17166 12189 17184 12223
rect 17132 12180 17184 12189
rect 17684 12180 17736 12232
rect 19156 12248 19208 12300
rect 23572 12359 23624 12368
rect 23572 12325 23581 12359
rect 23581 12325 23615 12359
rect 23615 12325 23624 12359
rect 23572 12316 23624 12325
rect 21364 12291 21416 12300
rect 21364 12257 21373 12291
rect 21373 12257 21407 12291
rect 21407 12257 21416 12291
rect 21364 12248 21416 12257
rect 21824 12291 21876 12300
rect 21824 12257 21833 12291
rect 21833 12257 21867 12291
rect 21867 12257 21876 12291
rect 21824 12248 21876 12257
rect 13268 12112 13320 12164
rect 15844 12112 15896 12164
rect 19800 12180 19852 12232
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 22100 12223 22152 12232
rect 22100 12189 22134 12223
rect 22134 12189 22152 12223
rect 22100 12180 22152 12189
rect 23204 12180 23256 12232
rect 22836 12112 22888 12164
rect 9404 12044 9456 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 13084 12044 13136 12096
rect 15292 12044 15344 12096
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 18604 12044 18656 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 19248 12044 19300 12096
rect 21088 12044 21140 12096
rect 21640 12044 21692 12096
rect 22192 12044 22244 12096
rect 2850 11942 2902 11994
rect 2914 11942 2966 11994
rect 2978 11942 3030 11994
rect 3042 11942 3094 11994
rect 3106 11942 3158 11994
rect 5850 11942 5902 11994
rect 5914 11942 5966 11994
rect 5978 11942 6030 11994
rect 6042 11942 6094 11994
rect 6106 11942 6158 11994
rect 8850 11942 8902 11994
rect 8914 11942 8966 11994
rect 8978 11942 9030 11994
rect 9042 11942 9094 11994
rect 9106 11942 9158 11994
rect 11850 11942 11902 11994
rect 11914 11942 11966 11994
rect 11978 11942 12030 11994
rect 12042 11942 12094 11994
rect 12106 11942 12158 11994
rect 14850 11942 14902 11994
rect 14914 11942 14966 11994
rect 14978 11942 15030 11994
rect 15042 11942 15094 11994
rect 15106 11942 15158 11994
rect 17850 11942 17902 11994
rect 17914 11942 17966 11994
rect 17978 11942 18030 11994
rect 18042 11942 18094 11994
rect 18106 11942 18158 11994
rect 20850 11942 20902 11994
rect 20914 11942 20966 11994
rect 20978 11942 21030 11994
rect 21042 11942 21094 11994
rect 21106 11942 21158 11994
rect 23850 11942 23902 11994
rect 23914 11942 23966 11994
rect 23978 11942 24030 11994
rect 24042 11942 24094 11994
rect 24106 11942 24158 11994
rect 388 11704 440 11756
rect 10876 11840 10928 11892
rect 11152 11840 11204 11892
rect 11704 11840 11756 11892
rect 3240 11704 3292 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 9220 11772 9272 11824
rect 9588 11772 9640 11824
rect 10692 11772 10744 11824
rect 14096 11840 14148 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 17684 11840 17736 11892
rect 18328 11840 18380 11892
rect 19248 11883 19300 11892
rect 19248 11849 19257 11883
rect 19257 11849 19291 11883
rect 19291 11849 19300 11883
rect 19248 11840 19300 11849
rect 9404 11747 9456 11756
rect 9404 11713 9438 11747
rect 9438 11713 9456 11747
rect 9404 11704 9456 11713
rect 10140 11704 10192 11756
rect 3332 11636 3384 11688
rect 4896 11636 4948 11688
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 7748 11636 7800 11688
rect 8484 11679 8536 11688
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 11060 11679 11112 11688
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 11152 11679 11204 11688
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 1676 11568 1728 11620
rect 11428 11568 11480 11620
rect 2780 11500 2832 11552
rect 3424 11500 3476 11552
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 8116 11543 8168 11552
rect 8116 11509 8125 11543
rect 8125 11509 8159 11543
rect 8159 11509 8168 11543
rect 8116 11500 8168 11509
rect 9404 11500 9456 11552
rect 13820 11772 13872 11824
rect 17408 11815 17460 11824
rect 17408 11781 17442 11815
rect 17442 11781 17460 11815
rect 17408 11772 17460 11781
rect 18696 11772 18748 11824
rect 21456 11840 21508 11892
rect 12716 11704 12768 11756
rect 12900 11704 12952 11756
rect 13084 11747 13136 11756
rect 13084 11713 13118 11747
rect 13118 11713 13136 11747
rect 13084 11704 13136 11713
rect 14188 11704 14240 11756
rect 16580 11704 16632 11756
rect 13728 11500 13780 11552
rect 15936 11568 15988 11620
rect 16856 11704 16908 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 23480 11772 23532 11824
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 23296 11747 23348 11756
rect 23296 11713 23305 11747
rect 23305 11713 23339 11747
rect 23339 11713 23348 11747
rect 23296 11704 23348 11713
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 21180 11636 21232 11688
rect 22836 11636 22888 11688
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 15660 11500 15712 11552
rect 16120 11500 16172 11552
rect 21272 11500 21324 11552
rect 21640 11543 21692 11552
rect 21640 11509 21649 11543
rect 21649 11509 21683 11543
rect 21683 11509 21692 11543
rect 21640 11500 21692 11509
rect 1350 11398 1402 11450
rect 1414 11398 1466 11450
rect 1478 11398 1530 11450
rect 1542 11398 1594 11450
rect 1606 11398 1658 11450
rect 4350 11398 4402 11450
rect 4414 11398 4466 11450
rect 4478 11398 4530 11450
rect 4542 11398 4594 11450
rect 4606 11398 4658 11450
rect 7350 11398 7402 11450
rect 7414 11398 7466 11450
rect 7478 11398 7530 11450
rect 7542 11398 7594 11450
rect 7606 11398 7658 11450
rect 10350 11398 10402 11450
rect 10414 11398 10466 11450
rect 10478 11398 10530 11450
rect 10542 11398 10594 11450
rect 10606 11398 10658 11450
rect 13350 11398 13402 11450
rect 13414 11398 13466 11450
rect 13478 11398 13530 11450
rect 13542 11398 13594 11450
rect 13606 11398 13658 11450
rect 16350 11398 16402 11450
rect 16414 11398 16466 11450
rect 16478 11398 16530 11450
rect 16542 11398 16594 11450
rect 16606 11398 16658 11450
rect 19350 11398 19402 11450
rect 19414 11398 19466 11450
rect 19478 11398 19530 11450
rect 19542 11398 19594 11450
rect 19606 11398 19658 11450
rect 22350 11398 22402 11450
rect 22414 11398 22466 11450
rect 22478 11398 22530 11450
rect 22542 11398 22594 11450
rect 22606 11398 22658 11450
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 8116 11296 8168 11348
rect 8668 11296 8720 11348
rect 11060 11296 11112 11348
rect 13084 11296 13136 11348
rect 13728 11296 13780 11348
rect 13820 11296 13872 11348
rect 16120 11296 16172 11348
rect 17500 11296 17552 11348
rect 3608 11271 3660 11280
rect 3608 11237 3617 11271
rect 3617 11237 3651 11271
rect 3651 11237 3660 11271
rect 3608 11228 3660 11237
rect 3516 11160 3568 11212
rect 3700 11160 3752 11212
rect 10692 11160 10744 11212
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 12532 11160 12584 11212
rect 12992 11160 13044 11212
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3792 11135 3844 11144
rect 3792 11101 3808 11135
rect 3808 11101 3842 11135
rect 3842 11101 3844 11135
rect 3792 11092 3844 11101
rect 5356 11092 5408 11144
rect 10140 11092 10192 11144
rect 14280 11160 14332 11212
rect 13268 11092 13320 11144
rect 15476 11228 15528 11280
rect 17316 11228 17368 11280
rect 18696 11296 18748 11348
rect 21824 11296 21876 11348
rect 20720 11228 20772 11280
rect 21456 11228 21508 11280
rect 3240 11024 3292 11076
rect 3608 11024 3660 11076
rect 6460 11024 6512 11076
rect 7012 11024 7064 11076
rect 8208 11024 8260 11076
rect 8944 11067 8996 11076
rect 8944 11033 8953 11067
rect 8953 11033 8987 11067
rect 8987 11033 8996 11067
rect 8944 11024 8996 11033
rect 9588 11024 9640 11076
rect 14004 11024 14056 11076
rect 14280 11067 14332 11076
rect 14280 11033 14289 11067
rect 14289 11033 14323 11067
rect 14323 11033 14332 11067
rect 14280 11024 14332 11033
rect 18328 11160 18380 11212
rect 21272 11160 21324 11212
rect 15660 11024 15712 11076
rect 16396 11067 16448 11076
rect 16396 11033 16405 11067
rect 16405 11033 16439 11067
rect 16439 11033 16448 11067
rect 16396 11024 16448 11033
rect 19800 11092 19852 11144
rect 20444 11092 20496 11144
rect 22008 11092 22060 11144
rect 20076 11024 20128 11076
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 3332 10956 3384 11008
rect 4252 10956 4304 11008
rect 5080 10956 5132 11008
rect 7748 10956 7800 11008
rect 8484 10956 8536 11008
rect 21272 10956 21324 11008
rect 23020 10956 23072 11008
rect 2850 10854 2902 10906
rect 2914 10854 2966 10906
rect 2978 10854 3030 10906
rect 3042 10854 3094 10906
rect 3106 10854 3158 10906
rect 5850 10854 5902 10906
rect 5914 10854 5966 10906
rect 5978 10854 6030 10906
rect 6042 10854 6094 10906
rect 6106 10854 6158 10906
rect 8850 10854 8902 10906
rect 8914 10854 8966 10906
rect 8978 10854 9030 10906
rect 9042 10854 9094 10906
rect 9106 10854 9158 10906
rect 11850 10854 11902 10906
rect 11914 10854 11966 10906
rect 11978 10854 12030 10906
rect 12042 10854 12094 10906
rect 12106 10854 12158 10906
rect 14850 10854 14902 10906
rect 14914 10854 14966 10906
rect 14978 10854 15030 10906
rect 15042 10854 15094 10906
rect 15106 10854 15158 10906
rect 17850 10854 17902 10906
rect 17914 10854 17966 10906
rect 17978 10854 18030 10906
rect 18042 10854 18094 10906
rect 18106 10854 18158 10906
rect 20850 10854 20902 10906
rect 20914 10854 20966 10906
rect 20978 10854 21030 10906
rect 21042 10854 21094 10906
rect 21106 10854 21158 10906
rect 23850 10854 23902 10906
rect 23914 10854 23966 10906
rect 23978 10854 24030 10906
rect 24042 10854 24094 10906
rect 24106 10854 24158 10906
rect 3332 10752 3384 10804
rect 2136 10684 2188 10736
rect 3424 10616 3476 10668
rect 5080 10752 5132 10804
rect 5448 10752 5500 10804
rect 7012 10752 7064 10804
rect 6184 10727 6236 10736
rect 6184 10693 6193 10727
rect 6193 10693 6227 10727
rect 6227 10693 6236 10727
rect 6184 10684 6236 10693
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 3516 10548 3568 10557
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 21180 10752 21232 10804
rect 21640 10752 21692 10804
rect 23388 10752 23440 10804
rect 11980 10684 12032 10736
rect 16396 10684 16448 10736
rect 21272 10727 21324 10736
rect 21272 10693 21281 10727
rect 21281 10693 21315 10727
rect 21315 10693 21324 10727
rect 21272 10684 21324 10693
rect 22008 10684 22060 10736
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7748 10616 7800 10668
rect 8484 10616 8536 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 11244 10616 11296 10668
rect 3884 10548 3936 10600
rect 4712 10548 4764 10600
rect 4896 10548 4948 10600
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 5632 10548 5684 10600
rect 8576 10548 8628 10600
rect 8760 10548 8812 10600
rect 9404 10548 9456 10600
rect 4068 10480 4120 10532
rect 7196 10480 7248 10532
rect 14096 10616 14148 10668
rect 19708 10659 19760 10668
rect 19708 10625 19742 10659
rect 19742 10625 19760 10659
rect 19708 10616 19760 10625
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 22100 10616 22152 10668
rect 15016 10548 15068 10600
rect 15844 10548 15896 10600
rect 12624 10480 12676 10532
rect 12992 10523 13044 10532
rect 12992 10489 13001 10523
rect 13001 10489 13035 10523
rect 13035 10489 13044 10523
rect 12992 10480 13044 10489
rect 1860 10412 1912 10464
rect 4896 10412 4948 10464
rect 6736 10412 6788 10464
rect 8300 10412 8352 10464
rect 8668 10412 8720 10464
rect 14464 10412 14516 10464
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16212 10412 16264 10464
rect 17316 10455 17368 10464
rect 17316 10421 17325 10455
rect 17325 10421 17359 10455
rect 17359 10421 17368 10455
rect 17316 10412 17368 10421
rect 21732 10548 21784 10600
rect 19800 10412 19852 10464
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 23572 10455 23624 10464
rect 23572 10421 23581 10455
rect 23581 10421 23615 10455
rect 23615 10421 23624 10455
rect 23572 10412 23624 10421
rect 1350 10310 1402 10362
rect 1414 10310 1466 10362
rect 1478 10310 1530 10362
rect 1542 10310 1594 10362
rect 1606 10310 1658 10362
rect 4350 10310 4402 10362
rect 4414 10310 4466 10362
rect 4478 10310 4530 10362
rect 4542 10310 4594 10362
rect 4606 10310 4658 10362
rect 7350 10310 7402 10362
rect 7414 10310 7466 10362
rect 7478 10310 7530 10362
rect 7542 10310 7594 10362
rect 7606 10310 7658 10362
rect 10350 10310 10402 10362
rect 10414 10310 10466 10362
rect 10478 10310 10530 10362
rect 10542 10310 10594 10362
rect 10606 10310 10658 10362
rect 13350 10310 13402 10362
rect 13414 10310 13466 10362
rect 13478 10310 13530 10362
rect 13542 10310 13594 10362
rect 13606 10310 13658 10362
rect 16350 10310 16402 10362
rect 16414 10310 16466 10362
rect 16478 10310 16530 10362
rect 16542 10310 16594 10362
rect 16606 10310 16658 10362
rect 19350 10310 19402 10362
rect 19414 10310 19466 10362
rect 19478 10310 19530 10362
rect 19542 10310 19594 10362
rect 19606 10310 19658 10362
rect 22350 10310 22402 10362
rect 22414 10310 22466 10362
rect 22478 10310 22530 10362
rect 22542 10310 22594 10362
rect 22606 10310 22658 10362
rect 4160 10208 4212 10260
rect 4804 10208 4856 10260
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 7748 10208 7800 10260
rect 8668 10208 8720 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 19708 10208 19760 10260
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 21272 10208 21324 10260
rect 3516 10140 3568 10192
rect 4160 10072 4212 10124
rect 12992 10140 13044 10192
rect 1768 9979 1820 9988
rect 1768 9945 1802 9979
rect 1802 9945 1820 9979
rect 1768 9936 1820 9945
rect 1860 9936 1912 9988
rect 3792 10004 3844 10056
rect 5356 10004 5408 10056
rect 6736 10047 6788 10056
rect 6736 10013 6754 10047
rect 6754 10013 6788 10047
rect 6736 10004 6788 10013
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 9588 10072 9640 10124
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 13728 10072 13780 10081
rect 15292 10183 15344 10192
rect 15292 10149 15301 10183
rect 15301 10149 15335 10183
rect 15335 10149 15344 10183
rect 15292 10140 15344 10149
rect 13176 10004 13228 10056
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 15844 10072 15896 10124
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 20904 10140 20956 10192
rect 23020 10251 23072 10260
rect 23020 10217 23029 10251
rect 23029 10217 23063 10251
rect 23063 10217 23072 10251
rect 23020 10208 23072 10217
rect 18512 10072 18564 10124
rect 4896 9979 4948 9988
rect 4896 9945 4914 9979
rect 4914 9945 4948 9979
rect 4896 9936 4948 9945
rect 3884 9868 3936 9920
rect 8300 9936 8352 9988
rect 8392 9936 8444 9988
rect 10508 9979 10560 9988
rect 10508 9945 10517 9979
rect 10517 9945 10551 9979
rect 10551 9945 10560 9979
rect 10508 9936 10560 9945
rect 11060 9936 11112 9988
rect 12440 9936 12492 9988
rect 14832 10004 14884 10056
rect 12532 9868 12584 9920
rect 13820 9868 13872 9920
rect 14188 9936 14240 9988
rect 16120 10004 16172 10056
rect 21180 10072 21232 10124
rect 21824 10072 21876 10124
rect 23572 10115 23624 10124
rect 23572 10081 23581 10115
rect 23581 10081 23615 10115
rect 23615 10081 23624 10115
rect 23572 10072 23624 10081
rect 20720 10004 20772 10056
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 22192 10004 22244 10056
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 16672 9979 16724 9988
rect 16672 9945 16706 9979
rect 16706 9945 16724 9979
rect 16672 9936 16724 9945
rect 16212 9911 16264 9920
rect 16212 9877 16221 9911
rect 16221 9877 16255 9911
rect 16255 9877 16264 9911
rect 16212 9868 16264 9877
rect 17132 9868 17184 9920
rect 22744 9868 22796 9920
rect 22836 9911 22888 9920
rect 22836 9877 22845 9911
rect 22845 9877 22879 9911
rect 22879 9877 22888 9911
rect 22836 9868 22888 9877
rect 2850 9766 2902 9818
rect 2914 9766 2966 9818
rect 2978 9766 3030 9818
rect 3042 9766 3094 9818
rect 3106 9766 3158 9818
rect 5850 9766 5902 9818
rect 5914 9766 5966 9818
rect 5978 9766 6030 9818
rect 6042 9766 6094 9818
rect 6106 9766 6158 9818
rect 8850 9766 8902 9818
rect 8914 9766 8966 9818
rect 8978 9766 9030 9818
rect 9042 9766 9094 9818
rect 9106 9766 9158 9818
rect 11850 9766 11902 9818
rect 11914 9766 11966 9818
rect 11978 9766 12030 9818
rect 12042 9766 12094 9818
rect 12106 9766 12158 9818
rect 14850 9766 14902 9818
rect 14914 9766 14966 9818
rect 14978 9766 15030 9818
rect 15042 9766 15094 9818
rect 15106 9766 15158 9818
rect 17850 9766 17902 9818
rect 17914 9766 17966 9818
rect 17978 9766 18030 9818
rect 18042 9766 18094 9818
rect 18106 9766 18158 9818
rect 20850 9766 20902 9818
rect 20914 9766 20966 9818
rect 20978 9766 21030 9818
rect 21042 9766 21094 9818
rect 21106 9766 21158 9818
rect 23850 9766 23902 9818
rect 23914 9766 23966 9818
rect 23978 9766 24030 9818
rect 24042 9766 24094 9818
rect 24106 9766 24158 9818
rect 1768 9664 1820 9716
rect 3240 9664 3292 9716
rect 3424 9664 3476 9716
rect 6368 9664 6420 9716
rect 7104 9664 7156 9716
rect 388 9528 440 9580
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 4160 9596 4212 9648
rect 2780 9392 2832 9444
rect 6644 9596 6696 9648
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 9312 9664 9364 9716
rect 10508 9707 10560 9716
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 14556 9664 14608 9716
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 8208 9639 8260 9648
rect 8208 9605 8217 9639
rect 8217 9605 8251 9639
rect 8251 9605 8260 9639
rect 8208 9596 8260 9605
rect 9220 9596 9272 9648
rect 15752 9707 15804 9716
rect 15752 9673 15761 9707
rect 15761 9673 15795 9707
rect 15795 9673 15804 9707
rect 15752 9664 15804 9673
rect 16672 9664 16724 9716
rect 17316 9664 17368 9716
rect 5264 9460 5316 9512
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 8392 9528 8444 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 6828 9460 6880 9512
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 9496 9460 9548 9512
rect 9680 9460 9732 9512
rect 12532 9528 12584 9580
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 14372 9571 14424 9580
rect 14372 9537 14381 9571
rect 14381 9537 14415 9571
rect 14415 9537 14424 9571
rect 14372 9528 14424 9537
rect 22652 9664 22704 9716
rect 14188 9460 14240 9512
rect 16764 9528 16816 9580
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 14556 9392 14608 9444
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 18236 9503 18288 9512
rect 16304 9392 16356 9444
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18420 9503 18472 9512
rect 18420 9469 18438 9503
rect 18438 9469 18472 9503
rect 18420 9460 18472 9469
rect 19800 9528 19852 9580
rect 6644 9324 6696 9376
rect 10784 9324 10836 9376
rect 12624 9324 12676 9376
rect 15292 9324 15344 9376
rect 19248 9503 19300 9512
rect 19248 9469 19257 9503
rect 19257 9469 19291 9503
rect 19291 9469 19300 9503
rect 19248 9460 19300 9469
rect 19064 9392 19116 9444
rect 19156 9392 19208 9444
rect 19616 9392 19668 9444
rect 20444 9392 20496 9444
rect 21272 9392 21324 9444
rect 18880 9324 18932 9376
rect 21180 9324 21232 9376
rect 21456 9571 21508 9580
rect 21456 9537 21465 9571
rect 21465 9537 21499 9571
rect 21499 9537 21508 9571
rect 21456 9528 21508 9537
rect 22008 9528 22060 9580
rect 22928 9528 22980 9580
rect 21548 9460 21600 9512
rect 22192 9392 22244 9444
rect 23388 9392 23440 9444
rect 22100 9324 22152 9376
rect 1350 9222 1402 9274
rect 1414 9222 1466 9274
rect 1478 9222 1530 9274
rect 1542 9222 1594 9274
rect 1606 9222 1658 9274
rect 4350 9222 4402 9274
rect 4414 9222 4466 9274
rect 4478 9222 4530 9274
rect 4542 9222 4594 9274
rect 4606 9222 4658 9274
rect 7350 9222 7402 9274
rect 7414 9222 7466 9274
rect 7478 9222 7530 9274
rect 7542 9222 7594 9274
rect 7606 9222 7658 9274
rect 10350 9222 10402 9274
rect 10414 9222 10466 9274
rect 10478 9222 10530 9274
rect 10542 9222 10594 9274
rect 10606 9222 10658 9274
rect 13350 9222 13402 9274
rect 13414 9222 13466 9274
rect 13478 9222 13530 9274
rect 13542 9222 13594 9274
rect 13606 9222 13658 9274
rect 16350 9222 16402 9274
rect 16414 9222 16466 9274
rect 16478 9222 16530 9274
rect 16542 9222 16594 9274
rect 16606 9222 16658 9274
rect 19350 9222 19402 9274
rect 19414 9222 19466 9274
rect 19478 9222 19530 9274
rect 19542 9222 19594 9274
rect 19606 9222 19658 9274
rect 22350 9222 22402 9274
rect 22414 9222 22466 9274
rect 22478 9222 22530 9274
rect 22542 9222 22594 9274
rect 22606 9222 22658 9274
rect 5816 9120 5868 9172
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 388 8916 440 8968
rect 2228 8823 2280 8832
rect 2228 8789 2237 8823
rect 2237 8789 2271 8823
rect 2271 8789 2280 8823
rect 2228 8780 2280 8789
rect 3700 9052 3752 9104
rect 5540 9052 5592 9104
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 5632 8984 5684 9036
rect 3240 8916 3292 8968
rect 4620 8916 4672 8968
rect 7932 8984 7984 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9588 8984 9640 9036
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 8668 8916 8720 8968
rect 11520 9120 11572 9172
rect 12440 9120 12492 9172
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 12900 9120 12952 9172
rect 15200 9120 15252 9172
rect 15844 9120 15896 9172
rect 16212 9120 16264 9172
rect 19156 9120 19208 9172
rect 19248 9120 19300 9172
rect 20720 9120 20772 9172
rect 22192 9120 22244 9172
rect 22928 9120 22980 9172
rect 19064 9052 19116 9104
rect 22008 9052 22060 9104
rect 15200 8984 15252 9036
rect 16028 9027 16080 9036
rect 16028 8993 16037 9027
rect 16037 8993 16071 9027
rect 16071 8993 16080 9027
rect 16028 8984 16080 8993
rect 23296 8984 23348 9036
rect 9496 8848 9548 8900
rect 12624 8916 12676 8968
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 16856 8916 16908 8968
rect 19800 8916 19852 8968
rect 21180 8959 21232 8968
rect 21180 8925 21214 8959
rect 21214 8925 21232 8959
rect 21180 8916 21232 8925
rect 22744 8916 22796 8968
rect 23388 8959 23440 8968
rect 23388 8925 23397 8959
rect 23397 8925 23431 8959
rect 23431 8925 23440 8959
rect 23388 8916 23440 8925
rect 11520 8848 11572 8900
rect 14740 8848 14792 8900
rect 16304 8891 16356 8900
rect 16304 8857 16338 8891
rect 16338 8857 16356 8891
rect 16304 8848 16356 8857
rect 17776 8891 17828 8900
rect 17776 8857 17810 8891
rect 17810 8857 17828 8891
rect 17776 8848 17828 8857
rect 18236 8848 18288 8900
rect 4160 8780 4212 8832
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 6368 8780 6420 8832
rect 8300 8780 8352 8832
rect 14648 8780 14700 8832
rect 16580 8780 16632 8832
rect 18420 8780 18472 8832
rect 19524 8891 19576 8900
rect 19524 8857 19558 8891
rect 19558 8857 19576 8891
rect 19524 8848 19576 8857
rect 21456 8848 21508 8900
rect 19892 8780 19944 8832
rect 2850 8678 2902 8730
rect 2914 8678 2966 8730
rect 2978 8678 3030 8730
rect 3042 8678 3094 8730
rect 3106 8678 3158 8730
rect 5850 8678 5902 8730
rect 5914 8678 5966 8730
rect 5978 8678 6030 8730
rect 6042 8678 6094 8730
rect 6106 8678 6158 8730
rect 8850 8678 8902 8730
rect 8914 8678 8966 8730
rect 8978 8678 9030 8730
rect 9042 8678 9094 8730
rect 9106 8678 9158 8730
rect 11850 8678 11902 8730
rect 11914 8678 11966 8730
rect 11978 8678 12030 8730
rect 12042 8678 12094 8730
rect 12106 8678 12158 8730
rect 14850 8678 14902 8730
rect 14914 8678 14966 8730
rect 14978 8678 15030 8730
rect 15042 8678 15094 8730
rect 15106 8678 15158 8730
rect 17850 8678 17902 8730
rect 17914 8678 17966 8730
rect 17978 8678 18030 8730
rect 18042 8678 18094 8730
rect 18106 8678 18158 8730
rect 20850 8678 20902 8730
rect 20914 8678 20966 8730
rect 20978 8678 21030 8730
rect 21042 8678 21094 8730
rect 21106 8678 21158 8730
rect 23850 8678 23902 8730
rect 23914 8678 23966 8730
rect 23978 8678 24030 8730
rect 24042 8678 24094 8730
rect 24106 8678 24158 8730
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 2228 8508 2280 8560
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 10140 8576 10192 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 14740 8576 14792 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 16764 8619 16816 8628
rect 16764 8585 16773 8619
rect 16773 8585 16807 8619
rect 16807 8585 16816 8619
rect 16764 8576 16816 8585
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 10048 8508 10100 8560
rect 15200 8508 15252 8560
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 19524 8576 19576 8628
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 1216 8304 1268 8356
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 4528 8372 4580 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 5724 8372 5776 8424
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 9220 8440 9272 8492
rect 9312 8372 9364 8424
rect 11704 8440 11756 8492
rect 14648 8440 14700 8492
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 18052 8551 18104 8560
rect 18052 8517 18061 8551
rect 18061 8517 18095 8551
rect 18095 8517 18104 8551
rect 18052 8508 18104 8517
rect 19800 8508 19852 8560
rect 14556 8372 14608 8424
rect 17868 8372 17920 8424
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 20628 8440 20680 8492
rect 20720 8440 20772 8492
rect 4896 8236 4948 8288
rect 16580 8304 16632 8356
rect 19892 8372 19944 8424
rect 20720 8304 20772 8356
rect 6920 8236 6972 8288
rect 9404 8236 9456 8288
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 17960 8236 18012 8288
rect 19708 8236 19760 8288
rect 1350 8134 1402 8186
rect 1414 8134 1466 8186
rect 1478 8134 1530 8186
rect 1542 8134 1594 8186
rect 1606 8134 1658 8186
rect 4350 8134 4402 8186
rect 4414 8134 4466 8186
rect 4478 8134 4530 8186
rect 4542 8134 4594 8186
rect 4606 8134 4658 8186
rect 7350 8134 7402 8186
rect 7414 8134 7466 8186
rect 7478 8134 7530 8186
rect 7542 8134 7594 8186
rect 7606 8134 7658 8186
rect 10350 8134 10402 8186
rect 10414 8134 10466 8186
rect 10478 8134 10530 8186
rect 10542 8134 10594 8186
rect 10606 8134 10658 8186
rect 13350 8134 13402 8186
rect 13414 8134 13466 8186
rect 13478 8134 13530 8186
rect 13542 8134 13594 8186
rect 13606 8134 13658 8186
rect 16350 8134 16402 8186
rect 16414 8134 16466 8186
rect 16478 8134 16530 8186
rect 16542 8134 16594 8186
rect 16606 8134 16658 8186
rect 19350 8134 19402 8186
rect 19414 8134 19466 8186
rect 19478 8134 19530 8186
rect 19542 8134 19594 8186
rect 19606 8134 19658 8186
rect 22350 8134 22402 8186
rect 22414 8134 22466 8186
rect 22478 8134 22530 8186
rect 22542 8134 22594 8186
rect 22606 8134 22658 8186
rect 3792 8032 3844 8084
rect 8024 8032 8076 8084
rect 4344 7964 4396 8016
rect 5724 8007 5776 8016
rect 5724 7973 5733 8007
rect 5733 7973 5767 8007
rect 5767 7973 5776 8007
rect 5724 7964 5776 7973
rect 7932 7964 7984 8016
rect 9220 8032 9272 8084
rect 13268 8032 13320 8084
rect 17776 8032 17828 8084
rect 19248 8075 19300 8084
rect 19248 8041 19257 8075
rect 19257 8041 19291 8075
rect 19291 8041 19300 8075
rect 19248 8032 19300 8041
rect 10140 7964 10192 8016
rect 12624 7964 12676 8016
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4160 7828 4212 7880
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 5540 7828 5592 7880
rect 3332 7760 3384 7812
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 4988 7760 5040 7812
rect 6920 7692 6972 7744
rect 8116 7896 8168 7948
rect 8852 7896 8904 7948
rect 7748 7760 7800 7812
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 9220 7828 9272 7880
rect 9496 7828 9548 7880
rect 11520 7828 11572 7880
rect 13176 7828 13228 7880
rect 17224 7964 17276 8016
rect 18052 7896 18104 7948
rect 18420 7939 18472 7948
rect 18420 7905 18429 7939
rect 18429 7905 18463 7939
rect 18463 7905 18472 7939
rect 18420 7896 18472 7905
rect 19708 7939 19760 7948
rect 19708 7905 19717 7939
rect 19717 7905 19751 7939
rect 19751 7905 19760 7939
rect 19708 7896 19760 7905
rect 19984 7896 20036 7948
rect 20720 8032 20772 8084
rect 21548 8032 21600 8084
rect 21824 7964 21876 8016
rect 20536 7896 20588 7948
rect 14004 7828 14056 7880
rect 14280 7828 14332 7880
rect 17960 7828 18012 7880
rect 19892 7828 19944 7880
rect 21272 7828 21324 7880
rect 8208 7760 8260 7812
rect 12716 7803 12768 7812
rect 12716 7769 12725 7803
rect 12725 7769 12759 7803
rect 12759 7769 12768 7803
rect 12716 7760 12768 7769
rect 9312 7692 9364 7744
rect 12256 7692 12308 7744
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 14556 7692 14608 7744
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 3042 7590 3094 7642
rect 3106 7590 3158 7642
rect 5850 7590 5902 7642
rect 5914 7590 5966 7642
rect 5978 7590 6030 7642
rect 6042 7590 6094 7642
rect 6106 7590 6158 7642
rect 8850 7590 8902 7642
rect 8914 7590 8966 7642
rect 8978 7590 9030 7642
rect 9042 7590 9094 7642
rect 9106 7590 9158 7642
rect 11850 7590 11902 7642
rect 11914 7590 11966 7642
rect 11978 7590 12030 7642
rect 12042 7590 12094 7642
rect 12106 7590 12158 7642
rect 14850 7590 14902 7642
rect 14914 7590 14966 7642
rect 14978 7590 15030 7642
rect 15042 7590 15094 7642
rect 15106 7590 15158 7642
rect 17850 7590 17902 7642
rect 17914 7590 17966 7642
rect 17978 7590 18030 7642
rect 18042 7590 18094 7642
rect 18106 7590 18158 7642
rect 20850 7590 20902 7642
rect 20914 7590 20966 7642
rect 20978 7590 21030 7642
rect 21042 7590 21094 7642
rect 21106 7590 21158 7642
rect 23850 7590 23902 7642
rect 23914 7590 23966 7642
rect 23978 7590 24030 7642
rect 24042 7590 24094 7642
rect 24106 7590 24158 7642
rect 3516 7488 3568 7540
rect 5540 7488 5592 7540
rect 8208 7488 8260 7540
rect 11704 7488 11756 7540
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 14280 7488 14332 7540
rect 19800 7488 19852 7540
rect 20536 7488 20588 7540
rect 20720 7488 20772 7540
rect 21548 7488 21600 7540
rect 3976 7420 4028 7472
rect 7196 7420 7248 7472
rect 4988 7352 5040 7404
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 6184 7284 6236 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8392 7352 8444 7404
rect 8484 7352 8536 7404
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9220 7352 9272 7404
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9588 7352 9640 7404
rect 12716 7420 12768 7472
rect 15200 7463 15252 7472
rect 15200 7429 15209 7463
rect 15209 7429 15243 7463
rect 15243 7429 15252 7463
rect 15200 7420 15252 7429
rect 12256 7352 12308 7404
rect 12440 7352 12492 7404
rect 8300 7284 8352 7336
rect 9496 7284 9548 7336
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 16856 7352 16908 7404
rect 17684 7352 17736 7404
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 20812 7352 20864 7404
rect 21364 7395 21416 7404
rect 21364 7361 21382 7395
rect 21382 7361 21416 7395
rect 21364 7352 21416 7361
rect 22836 7352 22888 7404
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 15476 7284 15528 7336
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 17960 7284 18012 7336
rect 15568 7216 15620 7268
rect 17776 7216 17828 7268
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 21640 7327 21692 7336
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 21732 7284 21784 7336
rect 4344 7148 4396 7200
rect 4712 7148 4764 7200
rect 8576 7148 8628 7200
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 16120 7148 16172 7200
rect 18420 7148 18472 7200
rect 18788 7148 18840 7200
rect 19708 7148 19760 7200
rect 23388 7148 23440 7200
rect 1350 7046 1402 7098
rect 1414 7046 1466 7098
rect 1478 7046 1530 7098
rect 1542 7046 1594 7098
rect 1606 7046 1658 7098
rect 4350 7046 4402 7098
rect 4414 7046 4466 7098
rect 4478 7046 4530 7098
rect 4542 7046 4594 7098
rect 4606 7046 4658 7098
rect 7350 7046 7402 7098
rect 7414 7046 7466 7098
rect 7478 7046 7530 7098
rect 7542 7046 7594 7098
rect 7606 7046 7658 7098
rect 10350 7046 10402 7098
rect 10414 7046 10466 7098
rect 10478 7046 10530 7098
rect 10542 7046 10594 7098
rect 10606 7046 10658 7098
rect 13350 7046 13402 7098
rect 13414 7046 13466 7098
rect 13478 7046 13530 7098
rect 13542 7046 13594 7098
rect 13606 7046 13658 7098
rect 16350 7046 16402 7098
rect 16414 7046 16466 7098
rect 16478 7046 16530 7098
rect 16542 7046 16594 7098
rect 16606 7046 16658 7098
rect 19350 7046 19402 7098
rect 19414 7046 19466 7098
rect 19478 7046 19530 7098
rect 19542 7046 19594 7098
rect 19606 7046 19658 7098
rect 22350 7046 22402 7098
rect 22414 7046 22466 7098
rect 22478 7046 22530 7098
rect 22542 7046 22594 7098
rect 22606 7046 22658 7098
rect 2872 6944 2924 6996
rect 7748 6944 7800 6996
rect 9128 6944 9180 6996
rect 12716 6944 12768 6996
rect 7840 6876 7892 6928
rect 4252 6808 4304 6860
rect 6920 6808 6972 6860
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 6184 6740 6236 6792
rect 7196 6672 7248 6724
rect 8024 6604 8076 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 8576 6672 8628 6724
rect 13268 6944 13320 6996
rect 20904 6944 20956 6996
rect 21732 6944 21784 6996
rect 13820 6876 13872 6928
rect 15568 6876 15620 6928
rect 20076 6876 20128 6928
rect 9220 6715 9272 6724
rect 9220 6681 9229 6715
rect 9229 6681 9263 6715
rect 9263 6681 9272 6715
rect 9220 6672 9272 6681
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 9772 6672 9824 6724
rect 9680 6604 9732 6656
rect 10048 6604 10100 6656
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 11704 6740 11756 6792
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 14464 6740 14516 6792
rect 15660 6808 15712 6860
rect 18880 6851 18932 6860
rect 18880 6817 18889 6851
rect 18889 6817 18923 6851
rect 18923 6817 18932 6851
rect 18880 6808 18932 6817
rect 19708 6808 19760 6860
rect 19800 6851 19852 6860
rect 19800 6817 19809 6851
rect 19809 6817 19843 6851
rect 19843 6817 19852 6851
rect 19800 6808 19852 6817
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 21456 6876 21508 6928
rect 20904 6808 20956 6860
rect 16764 6740 16816 6792
rect 17592 6740 17644 6792
rect 20168 6740 20220 6792
rect 12532 6672 12584 6724
rect 13176 6672 13228 6724
rect 12348 6604 12400 6656
rect 14004 6672 14056 6724
rect 15200 6672 15252 6724
rect 13820 6604 13872 6656
rect 15292 6604 15344 6656
rect 16028 6604 16080 6656
rect 16212 6604 16264 6656
rect 17960 6672 18012 6724
rect 18236 6672 18288 6724
rect 19064 6672 19116 6724
rect 19708 6672 19760 6724
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 21640 6740 21692 6792
rect 21824 6740 21876 6792
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 23112 6647 23164 6656
rect 23112 6613 23121 6647
rect 23121 6613 23155 6647
rect 23155 6613 23164 6647
rect 23112 6604 23164 6613
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 3042 6502 3094 6554
rect 3106 6502 3158 6554
rect 5850 6502 5902 6554
rect 5914 6502 5966 6554
rect 5978 6502 6030 6554
rect 6042 6502 6094 6554
rect 6106 6502 6158 6554
rect 8850 6502 8902 6554
rect 8914 6502 8966 6554
rect 8978 6502 9030 6554
rect 9042 6502 9094 6554
rect 9106 6502 9158 6554
rect 11850 6502 11902 6554
rect 11914 6502 11966 6554
rect 11978 6502 12030 6554
rect 12042 6502 12094 6554
rect 12106 6502 12158 6554
rect 14850 6502 14902 6554
rect 14914 6502 14966 6554
rect 14978 6502 15030 6554
rect 15042 6502 15094 6554
rect 15106 6502 15158 6554
rect 17850 6502 17902 6554
rect 17914 6502 17966 6554
rect 17978 6502 18030 6554
rect 18042 6502 18094 6554
rect 18106 6502 18158 6554
rect 20850 6502 20902 6554
rect 20914 6502 20966 6554
rect 20978 6502 21030 6554
rect 21042 6502 21094 6554
rect 21106 6502 21158 6554
rect 23850 6502 23902 6554
rect 23914 6502 23966 6554
rect 23978 6502 24030 6554
rect 24042 6502 24094 6554
rect 24106 6502 24158 6554
rect 8116 6400 8168 6452
rect 10140 6400 10192 6452
rect 11060 6400 11112 6452
rect 11612 6400 11664 6452
rect 11520 6332 11572 6384
rect 12256 6332 12308 6384
rect 9128 6264 9180 6316
rect 9312 6264 9364 6316
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 15752 6400 15804 6452
rect 17592 6400 17644 6452
rect 20076 6400 20128 6452
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 22836 6400 22888 6452
rect 14464 6332 14516 6384
rect 16028 6332 16080 6384
rect 18880 6332 18932 6384
rect 20168 6332 20220 6384
rect 9496 6264 9548 6273
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 14648 6264 14700 6316
rect 15200 6196 15252 6248
rect 18144 6264 18196 6316
rect 18512 6307 18564 6316
rect 18512 6273 18546 6307
rect 18546 6273 18564 6307
rect 18512 6264 18564 6273
rect 18972 6264 19024 6316
rect 21180 6307 21232 6316
rect 21180 6273 21189 6307
rect 21189 6273 21223 6307
rect 21223 6273 21232 6307
rect 21180 6264 21232 6273
rect 21640 6264 21692 6316
rect 23112 6332 23164 6384
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 19708 6239 19760 6248
rect 15476 6171 15528 6180
rect 15476 6137 15485 6171
rect 15485 6137 15519 6171
rect 15519 6137 15528 6171
rect 15476 6128 15528 6137
rect 16856 6128 16908 6180
rect 9680 6060 9732 6112
rect 13268 6103 13320 6112
rect 13268 6069 13277 6103
rect 13277 6069 13311 6103
rect 13311 6069 13320 6103
rect 13268 6060 13320 6069
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 16028 6060 16080 6112
rect 16948 6060 17000 6112
rect 17776 6060 17828 6112
rect 19708 6205 19717 6239
rect 19717 6205 19751 6239
rect 19751 6205 19760 6239
rect 19708 6196 19760 6205
rect 21548 6196 21600 6248
rect 21732 6128 21784 6180
rect 22192 6103 22244 6112
rect 22192 6069 22201 6103
rect 22201 6069 22235 6103
rect 22235 6069 22244 6103
rect 22192 6060 22244 6069
rect 1350 5958 1402 6010
rect 1414 5958 1466 6010
rect 1478 5958 1530 6010
rect 1542 5958 1594 6010
rect 1606 5958 1658 6010
rect 4350 5958 4402 6010
rect 4414 5958 4466 6010
rect 4478 5958 4530 6010
rect 4542 5958 4594 6010
rect 4606 5958 4658 6010
rect 7350 5958 7402 6010
rect 7414 5958 7466 6010
rect 7478 5958 7530 6010
rect 7542 5958 7594 6010
rect 7606 5958 7658 6010
rect 10350 5958 10402 6010
rect 10414 5958 10466 6010
rect 10478 5958 10530 6010
rect 10542 5958 10594 6010
rect 10606 5958 10658 6010
rect 13350 5958 13402 6010
rect 13414 5958 13466 6010
rect 13478 5958 13530 6010
rect 13542 5958 13594 6010
rect 13606 5958 13658 6010
rect 16350 5958 16402 6010
rect 16414 5958 16466 6010
rect 16478 5958 16530 6010
rect 16542 5958 16594 6010
rect 16606 5958 16658 6010
rect 19350 5958 19402 6010
rect 19414 5958 19466 6010
rect 19478 5958 19530 6010
rect 19542 5958 19594 6010
rect 19606 5958 19658 6010
rect 22350 5958 22402 6010
rect 22414 5958 22466 6010
rect 22478 5958 22530 6010
rect 22542 5958 22594 6010
rect 22606 5958 22658 6010
rect 9772 5899 9824 5908
rect 9772 5865 9781 5899
rect 9781 5865 9815 5899
rect 9815 5865 9824 5899
rect 9772 5856 9824 5865
rect 9864 5856 9916 5908
rect 12348 5856 12400 5908
rect 15476 5856 15528 5908
rect 5632 5720 5684 5772
rect 12440 5720 12492 5772
rect 14096 5763 14148 5772
rect 14096 5729 14105 5763
rect 14105 5729 14139 5763
rect 14139 5729 14148 5763
rect 14096 5720 14148 5729
rect 15476 5720 15528 5772
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 18972 5899 19024 5908
rect 18972 5865 18981 5899
rect 18981 5865 19015 5899
rect 19015 5865 19024 5899
rect 18972 5856 19024 5865
rect 19892 5856 19944 5908
rect 21272 5856 21324 5908
rect 16948 5788 17000 5840
rect 20444 5788 20496 5840
rect 18236 5720 18288 5772
rect 19708 5720 19760 5772
rect 22192 5788 22244 5840
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 6736 5584 6788 5636
rect 6828 5627 6880 5636
rect 6828 5593 6837 5627
rect 6837 5593 6871 5627
rect 6871 5593 6880 5627
rect 6828 5584 6880 5593
rect 7380 5652 7432 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 7196 5584 7248 5636
rect 8024 5584 8076 5636
rect 9680 5652 9732 5704
rect 9956 5652 10008 5704
rect 10048 5652 10100 5704
rect 14004 5652 14056 5704
rect 16304 5695 16356 5704
rect 16304 5661 16313 5695
rect 16313 5661 16347 5695
rect 16347 5661 16356 5695
rect 16304 5652 16356 5661
rect 17592 5652 17644 5704
rect 18328 5652 18380 5704
rect 18788 5695 18840 5704
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 21548 5652 21600 5704
rect 11520 5627 11572 5636
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 9404 5516 9456 5568
rect 12532 5584 12584 5636
rect 13268 5584 13320 5636
rect 20628 5584 20680 5636
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 17684 5516 17736 5568
rect 20720 5516 20772 5568
rect 21456 5516 21508 5568
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 3042 5414 3094 5466
rect 3106 5414 3158 5466
rect 5850 5414 5902 5466
rect 5914 5414 5966 5466
rect 5978 5414 6030 5466
rect 6042 5414 6094 5466
rect 6106 5414 6158 5466
rect 8850 5414 8902 5466
rect 8914 5414 8966 5466
rect 8978 5414 9030 5466
rect 9042 5414 9094 5466
rect 9106 5414 9158 5466
rect 11850 5414 11902 5466
rect 11914 5414 11966 5466
rect 11978 5414 12030 5466
rect 12042 5414 12094 5466
rect 12106 5414 12158 5466
rect 14850 5414 14902 5466
rect 14914 5414 14966 5466
rect 14978 5414 15030 5466
rect 15042 5414 15094 5466
rect 15106 5414 15158 5466
rect 17850 5414 17902 5466
rect 17914 5414 17966 5466
rect 17978 5414 18030 5466
rect 18042 5414 18094 5466
rect 18106 5414 18158 5466
rect 20850 5414 20902 5466
rect 20914 5414 20966 5466
rect 20978 5414 21030 5466
rect 21042 5414 21094 5466
rect 21106 5414 21158 5466
rect 23850 5414 23902 5466
rect 23914 5414 23966 5466
rect 23978 5414 24030 5466
rect 24042 5414 24094 5466
rect 24106 5414 24158 5466
rect 5632 5312 5684 5364
rect 6828 5312 6880 5364
rect 8668 5312 8720 5364
rect 8760 5312 8812 5364
rect 8944 5312 8996 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 15292 5312 15344 5321
rect 16212 5355 16264 5364
rect 16212 5321 16221 5355
rect 16221 5321 16255 5355
rect 16255 5321 16264 5355
rect 16212 5312 16264 5321
rect 16764 5312 16816 5364
rect 17500 5312 17552 5364
rect 6736 5244 6788 5296
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7380 5244 7432 5296
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7932 5244 7984 5296
rect 7748 5176 7800 5228
rect 8392 5244 8444 5296
rect 8852 5244 8904 5296
rect 8576 5176 8628 5228
rect 8668 5176 8720 5228
rect 15476 5176 15528 5228
rect 16120 5176 16172 5228
rect 16764 5176 16816 5228
rect 19984 5244 20036 5296
rect 7840 5108 7892 5160
rect 7196 5040 7248 5092
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 18236 5108 18288 5160
rect 20076 5219 20128 5228
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 8484 5040 8536 5092
rect 9404 5040 9456 5092
rect 19708 5040 19760 5092
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8024 4972 8076 5024
rect 12348 4972 12400 5024
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 21732 4972 21784 5024
rect 1350 4870 1402 4922
rect 1414 4870 1466 4922
rect 1478 4870 1530 4922
rect 1542 4870 1594 4922
rect 1606 4870 1658 4922
rect 4350 4870 4402 4922
rect 4414 4870 4466 4922
rect 4478 4870 4530 4922
rect 4542 4870 4594 4922
rect 4606 4870 4658 4922
rect 7350 4870 7402 4922
rect 7414 4870 7466 4922
rect 7478 4870 7530 4922
rect 7542 4870 7594 4922
rect 7606 4870 7658 4922
rect 10350 4870 10402 4922
rect 10414 4870 10466 4922
rect 10478 4870 10530 4922
rect 10542 4870 10594 4922
rect 10606 4870 10658 4922
rect 13350 4870 13402 4922
rect 13414 4870 13466 4922
rect 13478 4870 13530 4922
rect 13542 4870 13594 4922
rect 13606 4870 13658 4922
rect 16350 4870 16402 4922
rect 16414 4870 16466 4922
rect 16478 4870 16530 4922
rect 16542 4870 16594 4922
rect 16606 4870 16658 4922
rect 19350 4870 19402 4922
rect 19414 4870 19466 4922
rect 19478 4870 19530 4922
rect 19542 4870 19594 4922
rect 19606 4870 19658 4922
rect 22350 4870 22402 4922
rect 22414 4870 22466 4922
rect 22478 4870 22530 4922
rect 22542 4870 22594 4922
rect 22606 4870 22658 4922
rect 8208 4768 8260 4820
rect 5816 4632 5868 4684
rect 6920 4632 6972 4684
rect 7748 4700 7800 4752
rect 9220 4700 9272 4752
rect 9588 4700 9640 4752
rect 11520 4768 11572 4820
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 7840 4632 7892 4684
rect 6828 4564 6880 4616
rect 8668 4632 8720 4684
rect 8852 4632 8904 4684
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 18328 4632 18380 4684
rect 19800 4632 19852 4684
rect 20076 4632 20128 4684
rect 9588 4564 9640 4616
rect 7932 4496 7984 4548
rect 8576 4496 8628 4548
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 10968 4496 11020 4548
rect 16856 4496 16908 4548
rect 16948 4496 17000 4548
rect 5724 4428 5776 4480
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 7748 4428 7800 4480
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 9588 4471 9640 4480
rect 9588 4437 9597 4471
rect 9597 4437 9631 4471
rect 9631 4437 9640 4471
rect 9588 4428 9640 4437
rect 10784 4428 10836 4480
rect 12256 4428 12308 4480
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 19984 4564 20036 4616
rect 20260 4564 20312 4616
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 21272 4496 21324 4548
rect 17040 4428 17092 4437
rect 18880 4428 18932 4480
rect 19524 4428 19576 4480
rect 20076 4428 20128 4480
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 3042 4326 3094 4378
rect 3106 4326 3158 4378
rect 5850 4326 5902 4378
rect 5914 4326 5966 4378
rect 5978 4326 6030 4378
rect 6042 4326 6094 4378
rect 6106 4326 6158 4378
rect 8850 4326 8902 4378
rect 8914 4326 8966 4378
rect 8978 4326 9030 4378
rect 9042 4326 9094 4378
rect 9106 4326 9158 4378
rect 11850 4326 11902 4378
rect 11914 4326 11966 4378
rect 11978 4326 12030 4378
rect 12042 4326 12094 4378
rect 12106 4326 12158 4378
rect 14850 4326 14902 4378
rect 14914 4326 14966 4378
rect 14978 4326 15030 4378
rect 15042 4326 15094 4378
rect 15106 4326 15158 4378
rect 17850 4326 17902 4378
rect 17914 4326 17966 4378
rect 17978 4326 18030 4378
rect 18042 4326 18094 4378
rect 18106 4326 18158 4378
rect 20850 4326 20902 4378
rect 20914 4326 20966 4378
rect 20978 4326 21030 4378
rect 21042 4326 21094 4378
rect 21106 4326 21158 4378
rect 23850 4326 23902 4378
rect 23914 4326 23966 4378
rect 23978 4326 24030 4378
rect 24042 4326 24094 4378
rect 24106 4326 24158 4378
rect 6828 4224 6880 4276
rect 7288 4224 7340 4276
rect 9404 4224 9456 4276
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 17500 4224 17552 4276
rect 20352 4224 20404 4276
rect 21272 4267 21324 4276
rect 21272 4233 21281 4267
rect 21281 4233 21315 4267
rect 21315 4233 21324 4267
rect 21272 4224 21324 4233
rect 5724 4131 5776 4140
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 6276 4088 6328 4140
rect 6644 4088 6696 4140
rect 7932 4088 7984 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 6828 4020 6880 4072
rect 6920 4020 6972 4072
rect 8208 4020 8260 4072
rect 9404 4088 9456 4140
rect 10876 4156 10928 4208
rect 12256 4156 12308 4208
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 11704 4088 11756 4140
rect 13820 4156 13872 4208
rect 16212 4156 16264 4208
rect 13728 4131 13780 4140
rect 13728 4097 13762 4131
rect 13762 4097 13780 4131
rect 13728 4088 13780 4097
rect 15660 4088 15712 4140
rect 15936 4088 15988 4140
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 8300 3884 8352 3936
rect 9772 4020 9824 4072
rect 8760 3952 8812 4004
rect 9312 3952 9364 4004
rect 9864 3995 9916 4004
rect 9864 3961 9873 3995
rect 9873 3961 9907 3995
rect 9907 3961 9916 3995
rect 9864 3952 9916 3961
rect 10692 4020 10744 4072
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 14740 4020 14792 4072
rect 10876 3952 10928 4004
rect 16120 3952 16172 4004
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 9496 3884 9548 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 15384 3884 15436 3936
rect 15752 3884 15804 3936
rect 17132 4088 17184 4140
rect 17408 4088 17460 4140
rect 18328 4088 18380 4140
rect 19708 4088 19760 4140
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 20352 4131 20404 4140
rect 20352 4097 20386 4131
rect 20386 4097 20404 4131
rect 20352 4088 20404 4097
rect 21456 4131 21508 4140
rect 21456 4097 21465 4131
rect 21465 4097 21499 4131
rect 21499 4097 21508 4131
rect 21456 4088 21508 4097
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 17776 4063 17828 4072
rect 17776 4029 17785 4063
rect 17785 4029 17819 4063
rect 17819 4029 17828 4063
rect 17776 4020 17828 4029
rect 19524 4063 19576 4072
rect 19524 4029 19533 4063
rect 19533 4029 19567 4063
rect 19567 4029 19576 4063
rect 19524 4020 19576 4029
rect 16856 3952 16908 4004
rect 20720 4020 20772 4072
rect 19892 3952 19944 4004
rect 20076 3884 20128 3936
rect 21640 3884 21692 3936
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 1350 3782 1402 3834
rect 1414 3782 1466 3834
rect 1478 3782 1530 3834
rect 1542 3782 1594 3834
rect 1606 3782 1658 3834
rect 4350 3782 4402 3834
rect 4414 3782 4466 3834
rect 4478 3782 4530 3834
rect 4542 3782 4594 3834
rect 4606 3782 4658 3834
rect 7350 3782 7402 3834
rect 7414 3782 7466 3834
rect 7478 3782 7530 3834
rect 7542 3782 7594 3834
rect 7606 3782 7658 3834
rect 10350 3782 10402 3834
rect 10414 3782 10466 3834
rect 10478 3782 10530 3834
rect 10542 3782 10594 3834
rect 10606 3782 10658 3834
rect 13350 3782 13402 3834
rect 13414 3782 13466 3834
rect 13478 3782 13530 3834
rect 13542 3782 13594 3834
rect 13606 3782 13658 3834
rect 16350 3782 16402 3834
rect 16414 3782 16466 3834
rect 16478 3782 16530 3834
rect 16542 3782 16594 3834
rect 16606 3782 16658 3834
rect 19350 3782 19402 3834
rect 19414 3782 19466 3834
rect 19478 3782 19530 3834
rect 19542 3782 19594 3834
rect 19606 3782 19658 3834
rect 22350 3782 22402 3834
rect 22414 3782 22466 3834
rect 22478 3782 22530 3834
rect 22542 3782 22594 3834
rect 22606 3782 22658 3834
rect 8392 3680 8444 3732
rect 9036 3680 9088 3732
rect 9220 3680 9272 3732
rect 10232 3680 10284 3732
rect 10784 3680 10836 3732
rect 13728 3680 13780 3732
rect 16028 3680 16080 3732
rect 4712 3544 4764 3596
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 7932 3612 7984 3664
rect 8024 3655 8076 3664
rect 8024 3621 8033 3655
rect 8033 3621 8067 3655
rect 8067 3621 8076 3655
rect 8024 3612 8076 3621
rect 8668 3612 8720 3664
rect 9496 3655 9548 3664
rect 6828 3544 6880 3596
rect 8300 3544 8352 3596
rect 8484 3544 8536 3596
rect 9496 3621 9505 3655
rect 9505 3621 9539 3655
rect 9539 3621 9548 3655
rect 9496 3612 9548 3621
rect 9772 3612 9824 3664
rect 7748 3476 7800 3528
rect 7288 3408 7340 3460
rect 8392 3476 8444 3528
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 10784 3544 10836 3596
rect 13820 3544 13872 3596
rect 9588 3476 9640 3528
rect 14648 3544 14700 3596
rect 16120 3587 16172 3596
rect 16120 3553 16138 3587
rect 16138 3553 16172 3587
rect 16120 3544 16172 3553
rect 17040 3544 17092 3596
rect 18236 3680 18288 3732
rect 19708 3680 19760 3732
rect 20444 3680 20496 3732
rect 14924 3476 14976 3528
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15292 3476 15344 3528
rect 15936 3519 15988 3528
rect 15936 3485 15945 3519
rect 15945 3485 15979 3519
rect 15979 3485 15988 3519
rect 15936 3476 15988 3485
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 17776 3476 17828 3528
rect 9036 3408 9088 3460
rect 9496 3408 9548 3460
rect 9864 3451 9916 3460
rect 9864 3417 9873 3451
rect 9873 3417 9907 3451
rect 9907 3417 9916 3451
rect 9864 3408 9916 3417
rect 7564 3340 7616 3392
rect 8300 3340 8352 3392
rect 9404 3340 9456 3392
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 10232 3408 10284 3460
rect 12164 3408 12216 3460
rect 13176 3451 13228 3460
rect 13176 3417 13185 3451
rect 13185 3417 13219 3451
rect 13219 3417 13228 3451
rect 13176 3408 13228 3417
rect 17316 3408 17368 3460
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 21364 3476 21416 3528
rect 21640 3544 21692 3596
rect 21732 3476 21784 3528
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 10876 3340 10928 3349
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 17132 3340 17184 3392
rect 18696 3383 18748 3392
rect 18696 3349 18705 3383
rect 18705 3349 18739 3383
rect 18739 3349 18748 3383
rect 18696 3340 18748 3349
rect 19708 3340 19760 3392
rect 21916 3383 21968 3392
rect 21916 3349 21925 3383
rect 21925 3349 21959 3383
rect 21959 3349 21968 3383
rect 21916 3340 21968 3349
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 3042 3238 3094 3290
rect 3106 3238 3158 3290
rect 5850 3238 5902 3290
rect 5914 3238 5966 3290
rect 5978 3238 6030 3290
rect 6042 3238 6094 3290
rect 6106 3238 6158 3290
rect 8850 3238 8902 3290
rect 8914 3238 8966 3290
rect 8978 3238 9030 3290
rect 9042 3238 9094 3290
rect 9106 3238 9158 3290
rect 11850 3238 11902 3290
rect 11914 3238 11966 3290
rect 11978 3238 12030 3290
rect 12042 3238 12094 3290
rect 12106 3238 12158 3290
rect 14850 3238 14902 3290
rect 14914 3238 14966 3290
rect 14978 3238 15030 3290
rect 15042 3238 15094 3290
rect 15106 3238 15158 3290
rect 17850 3238 17902 3290
rect 17914 3238 17966 3290
rect 17978 3238 18030 3290
rect 18042 3238 18094 3290
rect 18106 3238 18158 3290
rect 20850 3238 20902 3290
rect 20914 3238 20966 3290
rect 20978 3238 21030 3290
rect 21042 3238 21094 3290
rect 21106 3238 21158 3290
rect 23850 3238 23902 3290
rect 23914 3238 23966 3290
rect 23978 3238 24030 3290
rect 24042 3238 24094 3290
rect 24106 3238 24158 3290
rect 7564 3136 7616 3188
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 9496 3136 9548 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 7932 3068 7984 3120
rect 8208 3068 8260 3120
rect 11336 3136 11388 3188
rect 13176 3136 13228 3188
rect 14740 3136 14792 3188
rect 15200 3136 15252 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 10692 3111 10744 3120
rect 10692 3077 10701 3111
rect 10701 3077 10735 3111
rect 10735 3077 10744 3111
rect 10692 3068 10744 3077
rect 6184 3000 6236 3052
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10048 3000 10100 3052
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 13820 3068 13872 3120
rect 15292 3111 15344 3120
rect 15292 3077 15301 3111
rect 15301 3077 15335 3111
rect 15335 3077 15344 3111
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 19708 3179 19760 3188
rect 19708 3145 19717 3179
rect 19717 3145 19751 3179
rect 19751 3145 19760 3179
rect 19708 3136 19760 3145
rect 21456 3136 21508 3188
rect 15292 3068 15344 3077
rect 9588 2932 9640 2984
rect 10232 2932 10284 2984
rect 9496 2864 9548 2916
rect 13728 3043 13780 3052
rect 13728 3009 13762 3043
rect 13762 3009 13780 3043
rect 13728 3000 13780 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 17316 3068 17368 3120
rect 18696 3068 18748 3120
rect 19800 3068 19852 3120
rect 21824 3068 21876 3120
rect 17040 3000 17092 3052
rect 17132 3000 17184 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 15568 2975 15620 2984
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 17224 2932 17276 2984
rect 20628 3000 20680 3052
rect 7288 2796 7340 2848
rect 10140 2796 10192 2848
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 19984 2864 20036 2916
rect 19248 2839 19300 2848
rect 19248 2805 19257 2839
rect 19257 2805 19291 2839
rect 19291 2805 19300 2839
rect 19248 2796 19300 2805
rect 1350 2694 1402 2746
rect 1414 2694 1466 2746
rect 1478 2694 1530 2746
rect 1542 2694 1594 2746
rect 1606 2694 1658 2746
rect 4350 2694 4402 2746
rect 4414 2694 4466 2746
rect 4478 2694 4530 2746
rect 4542 2694 4594 2746
rect 4606 2694 4658 2746
rect 7350 2694 7402 2746
rect 7414 2694 7466 2746
rect 7478 2694 7530 2746
rect 7542 2694 7594 2746
rect 7606 2694 7658 2746
rect 10350 2694 10402 2746
rect 10414 2694 10466 2746
rect 10478 2694 10530 2746
rect 10542 2694 10594 2746
rect 10606 2694 10658 2746
rect 13350 2694 13402 2746
rect 13414 2694 13466 2746
rect 13478 2694 13530 2746
rect 13542 2694 13594 2746
rect 13606 2694 13658 2746
rect 16350 2694 16402 2746
rect 16414 2694 16466 2746
rect 16478 2694 16530 2746
rect 16542 2694 16594 2746
rect 16606 2694 16658 2746
rect 19350 2694 19402 2746
rect 19414 2694 19466 2746
rect 19478 2694 19530 2746
rect 19542 2694 19594 2746
rect 19606 2694 19658 2746
rect 22350 2694 22402 2746
rect 22414 2694 22466 2746
rect 22478 2694 22530 2746
rect 22542 2694 22594 2746
rect 22606 2694 22658 2746
rect 7196 2592 7248 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 12992 2592 13044 2644
rect 14372 2592 14424 2644
rect 15292 2592 15344 2644
rect 16764 2592 16816 2644
rect 18328 2592 18380 2644
rect 19708 2592 19760 2644
rect 8024 2524 8076 2576
rect 5724 2388 5776 2440
rect 6736 2388 6788 2440
rect 8300 2456 8352 2508
rect 12532 2524 12584 2576
rect 9680 2456 9732 2508
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 8576 2388 8628 2440
rect 9220 2388 9272 2440
rect 7104 2320 7156 2372
rect 7748 2363 7800 2372
rect 7748 2329 7757 2363
rect 7757 2329 7791 2363
rect 7791 2329 7800 2363
rect 7748 2320 7800 2329
rect 9680 2320 9732 2372
rect 17500 2456 17552 2508
rect 10324 2388 10376 2440
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 11612 2388 11664 2440
rect 12808 2388 12860 2440
rect 14188 2388 14240 2440
rect 14556 2388 14608 2440
rect 15476 2388 15528 2440
rect 16120 2388 16172 2440
rect 19248 2388 19300 2440
rect 19340 2388 19392 2440
rect 21916 2431 21968 2440
rect 21916 2397 21925 2431
rect 21925 2397 21959 2431
rect 21959 2397 21968 2431
rect 21916 2388 21968 2397
rect 12256 2320 12308 2372
rect 16764 2320 16816 2372
rect 17408 2320 17460 2372
rect 18420 2320 18472 2372
rect 6460 2252 6512 2304
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 14740 2252 14792 2304
rect 21272 2252 21324 2304
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 3042 2150 3094 2202
rect 3106 2150 3158 2202
rect 5850 2150 5902 2202
rect 5914 2150 5966 2202
rect 5978 2150 6030 2202
rect 6042 2150 6094 2202
rect 6106 2150 6158 2202
rect 8850 2150 8902 2202
rect 8914 2150 8966 2202
rect 8978 2150 9030 2202
rect 9042 2150 9094 2202
rect 9106 2150 9158 2202
rect 11850 2150 11902 2202
rect 11914 2150 11966 2202
rect 11978 2150 12030 2202
rect 12042 2150 12094 2202
rect 12106 2150 12158 2202
rect 14850 2150 14902 2202
rect 14914 2150 14966 2202
rect 14978 2150 15030 2202
rect 15042 2150 15094 2202
rect 15106 2150 15158 2202
rect 17850 2150 17902 2202
rect 17914 2150 17966 2202
rect 17978 2150 18030 2202
rect 18042 2150 18094 2202
rect 18106 2150 18158 2202
rect 20850 2150 20902 2202
rect 20914 2150 20966 2202
rect 20978 2150 21030 2202
rect 21042 2150 21094 2202
rect 21106 2150 21158 2202
rect 23850 2150 23902 2202
rect 23914 2150 23966 2202
rect 23978 2150 24030 2202
rect 24042 2150 24094 2202
rect 24106 2150 24158 2202
<< metal2 >>
rect 5170 26924 5226 27324
rect 5552 26982 5764 27010
rect 2850 25052 3158 25061
rect 2850 25050 2856 25052
rect 2912 25050 2936 25052
rect 2992 25050 3016 25052
rect 3072 25050 3096 25052
rect 3152 25050 3158 25052
rect 2912 24998 2914 25050
rect 3094 24998 3096 25050
rect 2850 24996 2856 24998
rect 2912 24996 2936 24998
rect 2992 24996 3016 24998
rect 3072 24996 3096 24998
rect 3152 24996 3158 24998
rect 2850 24987 3158 24996
rect 5184 24818 5212 26924
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 5172 24676 5224 24682
rect 5172 24618 5224 24624
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 1350 24508 1658 24517
rect 1350 24506 1356 24508
rect 1412 24506 1436 24508
rect 1492 24506 1516 24508
rect 1572 24506 1596 24508
rect 1652 24506 1658 24508
rect 1412 24454 1414 24506
rect 1594 24454 1596 24506
rect 1350 24452 1356 24454
rect 1412 24452 1436 24454
rect 1492 24452 1516 24454
rect 1572 24452 1596 24454
rect 1652 24452 1658 24454
rect 1350 24443 1658 24452
rect 4350 24508 4658 24517
rect 4350 24506 4356 24508
rect 4412 24506 4436 24508
rect 4492 24506 4516 24508
rect 4572 24506 4596 24508
rect 4652 24506 4658 24508
rect 4412 24454 4414 24506
rect 4594 24454 4596 24506
rect 4350 24452 4356 24454
rect 4412 24452 4436 24454
rect 4492 24452 4516 24454
rect 4572 24452 4596 24454
rect 4652 24452 4658 24454
rect 4350 24443 4658 24452
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 2850 23964 3158 23973
rect 2850 23962 2856 23964
rect 2912 23962 2936 23964
rect 2992 23962 3016 23964
rect 3072 23962 3096 23964
rect 3152 23962 3158 23964
rect 2912 23910 2914 23962
rect 3094 23910 3096 23962
rect 2850 23908 2856 23910
rect 2912 23908 2936 23910
rect 2992 23908 3016 23910
rect 3072 23908 3096 23910
rect 3152 23908 3158 23910
rect 2850 23899 3158 23908
rect 3436 23866 3464 24074
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3528 23730 3556 24142
rect 4252 23792 4304 23798
rect 4252 23734 4304 23740
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 1350 23420 1658 23429
rect 1350 23418 1356 23420
rect 1412 23418 1436 23420
rect 1492 23418 1516 23420
rect 1572 23418 1596 23420
rect 1652 23418 1658 23420
rect 1412 23366 1414 23418
rect 1594 23366 1596 23418
rect 1350 23364 1356 23366
rect 1412 23364 1436 23366
rect 1492 23364 1516 23366
rect 1572 23364 1596 23366
rect 1652 23364 1658 23366
rect 1350 23355 1658 23364
rect 3804 23322 3832 23666
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 2850 22876 3158 22885
rect 2850 22874 2856 22876
rect 2912 22874 2936 22876
rect 2992 22874 3016 22876
rect 3072 22874 3096 22876
rect 3152 22874 3158 22876
rect 2912 22822 2914 22874
rect 3094 22822 3096 22874
rect 2850 22820 2856 22822
rect 2912 22820 2936 22822
rect 2992 22820 3016 22822
rect 3072 22820 3096 22822
rect 3152 22820 3158 22822
rect 2850 22811 3158 22820
rect 4264 22778 4292 23734
rect 4350 23420 4658 23429
rect 4350 23418 4356 23420
rect 4412 23418 4436 23420
rect 4492 23418 4516 23420
rect 4572 23418 4596 23420
rect 4652 23418 4658 23420
rect 4412 23366 4414 23418
rect 4594 23366 4596 23418
rect 4350 23364 4356 23366
rect 4412 23364 4436 23366
rect 4492 23364 4516 23366
rect 4572 23364 4596 23366
rect 4652 23364 4658 23366
rect 4350 23355 4658 23364
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4724 22778 4752 22918
rect 4252 22772 4304 22778
rect 4252 22714 4304 22720
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4816 22710 4844 22918
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 5000 22642 5028 24550
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 1350 22332 1658 22341
rect 1350 22330 1356 22332
rect 1412 22330 1436 22332
rect 1492 22330 1516 22332
rect 1572 22330 1596 22332
rect 1652 22330 1658 22332
rect 1412 22278 1414 22330
rect 1594 22278 1596 22330
rect 1350 22276 1356 22278
rect 1412 22276 1436 22278
rect 1492 22276 1516 22278
rect 1572 22276 1596 22278
rect 1652 22276 1658 22278
rect 1350 22267 1658 22276
rect 4350 22332 4658 22341
rect 4350 22330 4356 22332
rect 4412 22330 4436 22332
rect 4492 22330 4516 22332
rect 4572 22330 4596 22332
rect 4652 22330 4658 22332
rect 4412 22278 4414 22330
rect 4594 22278 4596 22330
rect 4350 22276 4356 22278
rect 4412 22276 4436 22278
rect 4492 22276 4516 22278
rect 4572 22276 4596 22278
rect 4652 22276 4658 22278
rect 4350 22267 4658 22276
rect 4908 22234 4936 22510
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 2850 21788 3158 21797
rect 2850 21786 2856 21788
rect 2912 21786 2936 21788
rect 2992 21786 3016 21788
rect 3072 21786 3096 21788
rect 3152 21786 3158 21788
rect 2912 21734 2914 21786
rect 3094 21734 3096 21786
rect 2850 21732 2856 21734
rect 2912 21732 2936 21734
rect 2992 21732 3016 21734
rect 3072 21732 3096 21734
rect 3152 21732 3158 21734
rect 2850 21723 3158 21732
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 1350 21244 1658 21253
rect 1350 21242 1356 21244
rect 1412 21242 1436 21244
rect 1492 21242 1516 21244
rect 1572 21242 1596 21244
rect 1652 21242 1658 21244
rect 1412 21190 1414 21242
rect 1594 21190 1596 21242
rect 1350 21188 1356 21190
rect 1412 21188 1436 21190
rect 1492 21188 1516 21190
rect 1572 21188 1596 21190
rect 1652 21188 1658 21190
rect 1350 21179 1658 21188
rect 3804 21146 3832 21490
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 2850 20700 3158 20709
rect 2850 20698 2856 20700
rect 2912 20698 2936 20700
rect 2992 20698 3016 20700
rect 3072 20698 3096 20700
rect 3152 20698 3158 20700
rect 2912 20646 2914 20698
rect 3094 20646 3096 20698
rect 2850 20644 2856 20646
rect 2912 20644 2936 20646
rect 2992 20644 3016 20646
rect 3072 20644 3096 20646
rect 3152 20644 3158 20646
rect 2850 20635 3158 20644
rect 3528 20466 3556 20742
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 4172 20262 4200 21286
rect 4264 20942 4292 21830
rect 4632 21350 4660 21966
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4350 21244 4658 21253
rect 4350 21242 4356 21244
rect 4412 21242 4436 21244
rect 4492 21242 4516 21244
rect 4572 21242 4596 21244
rect 4652 21242 4658 21244
rect 4412 21190 4414 21242
rect 4594 21190 4596 21242
rect 4350 21188 4356 21190
rect 4412 21188 4436 21190
rect 4492 21188 4516 21190
rect 4572 21188 4596 21190
rect 4652 21188 4658 21190
rect 4350 21179 4658 21188
rect 4724 21146 4752 21830
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 4816 20942 4844 21898
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 5092 20466 5120 22374
rect 5184 22098 5212 24618
rect 5552 24206 5580 26982
rect 5736 26874 5764 26982
rect 5814 26924 5870 27324
rect 6458 26924 6514 27324
rect 7102 26924 7158 27324
rect 8390 26924 8446 27324
rect 8772 26982 8984 27010
rect 5828 26874 5856 26924
rect 5736 26846 5856 26874
rect 5850 25052 6158 25061
rect 5850 25050 5856 25052
rect 5912 25050 5936 25052
rect 5992 25050 6016 25052
rect 6072 25050 6096 25052
rect 6152 25050 6158 25052
rect 5912 24998 5914 25050
rect 6094 24998 6096 25050
rect 5850 24996 5856 24998
rect 5912 24996 5936 24998
rect 5992 24996 6016 24998
rect 6072 24996 6096 24998
rect 6152 24996 6158 24998
rect 5850 24987 6158 24996
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5644 24342 5672 24686
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5632 24336 5684 24342
rect 5632 24278 5684 24284
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 5460 23866 5488 24006
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5644 23746 5672 24278
rect 5736 23866 5764 24618
rect 6472 24614 6500 26924
rect 6552 24744 6604 24750
rect 6552 24686 6604 24692
rect 6460 24608 6512 24614
rect 6460 24550 6512 24556
rect 5850 23964 6158 23973
rect 5850 23962 5856 23964
rect 5912 23962 5936 23964
rect 5992 23962 6016 23964
rect 6072 23962 6096 23964
rect 6152 23962 6158 23964
rect 5912 23910 5914 23962
rect 6094 23910 6096 23962
rect 5850 23908 5856 23910
rect 5912 23908 5936 23910
rect 5992 23908 6016 23910
rect 6072 23908 6096 23910
rect 6152 23908 6158 23910
rect 5850 23899 6158 23908
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5644 23718 5764 23746
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5448 23180 5500 23186
rect 5500 23140 5580 23168
rect 5448 23122 5500 23128
rect 5276 22710 5304 23122
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5170 21992 5226 22001
rect 5170 21927 5226 21936
rect 5184 21622 5212 21927
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5276 21010 5304 22646
rect 5552 22114 5580 23140
rect 5644 22642 5672 23462
rect 5736 23168 5764 23718
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 6104 23186 6132 23462
rect 5908 23180 5960 23186
rect 5736 23140 5908 23168
rect 5908 23122 5960 23128
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 5850 22876 6158 22885
rect 5850 22874 5856 22876
rect 5912 22874 5936 22876
rect 5992 22874 6016 22876
rect 6072 22874 6096 22876
rect 6152 22874 6158 22876
rect 5912 22822 5914 22874
rect 6094 22822 6096 22874
rect 5850 22820 5856 22822
rect 5912 22820 5936 22822
rect 5992 22820 6016 22822
rect 6072 22820 6096 22822
rect 6152 22820 6158 22822
rect 5850 22811 6158 22820
rect 6288 22778 6316 23598
rect 6564 23594 6592 24686
rect 7116 24614 7144 26924
rect 8404 24818 8432 26924
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6748 23730 6776 24346
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 6552 23588 6604 23594
rect 6552 23530 6604 23536
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 5552 22086 5764 22114
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 1350 20156 1658 20165
rect 1350 20154 1356 20156
rect 1412 20154 1436 20156
rect 1492 20154 1516 20156
rect 1572 20154 1596 20156
rect 1652 20154 1658 20156
rect 1412 20102 1414 20154
rect 1594 20102 1596 20154
rect 1350 20100 1356 20102
rect 1412 20100 1436 20102
rect 1492 20100 1516 20102
rect 1572 20100 1596 20102
rect 1652 20100 1658 20102
rect 1350 20091 1658 20100
rect 2850 19612 3158 19621
rect 2850 19610 2856 19612
rect 2912 19610 2936 19612
rect 2992 19610 3016 19612
rect 3072 19610 3096 19612
rect 3152 19610 3158 19612
rect 2912 19558 2914 19610
rect 3094 19558 3096 19610
rect 2850 19556 2856 19558
rect 2912 19556 2936 19558
rect 2992 19556 3016 19558
rect 3072 19556 3096 19558
rect 3152 19556 3158 19558
rect 2850 19547 3158 19556
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 1216 19168 1268 19174
rect 1214 19136 1216 19145
rect 1268 19136 1270 19145
rect 1214 19071 1270 19080
rect 1350 19068 1658 19077
rect 1350 19066 1356 19068
rect 1412 19066 1436 19068
rect 1492 19066 1516 19068
rect 1572 19066 1596 19068
rect 1652 19066 1658 19068
rect 1412 19014 1414 19066
rect 1594 19014 1596 19066
rect 1350 19012 1356 19014
rect 1412 19012 1436 19014
rect 1492 19012 1516 19014
rect 1572 19012 1596 19014
rect 1652 19012 1658 19014
rect 1350 19003 1658 19012
rect 3528 18970 3556 19314
rect 4172 19174 4200 20198
rect 4350 20156 4658 20165
rect 4350 20154 4356 20156
rect 4412 20154 4436 20156
rect 4492 20154 4516 20156
rect 4572 20154 4596 20156
rect 4652 20154 4658 20156
rect 4412 20102 4414 20154
rect 4594 20102 4596 20154
rect 4350 20100 4356 20102
rect 4412 20100 4436 20102
rect 4492 20100 4516 20102
rect 4572 20100 4596 20102
rect 4652 20100 4658 20102
rect 4350 20091 4658 20100
rect 5276 19530 5304 20946
rect 5460 20534 5488 21422
rect 5644 21010 5672 21966
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5644 20602 5672 20946
rect 5736 20924 5764 22086
rect 5850 21788 6158 21797
rect 5850 21786 5856 21788
rect 5912 21786 5936 21788
rect 5992 21786 6016 21788
rect 6072 21786 6096 21788
rect 6152 21786 6158 21788
rect 5912 21734 5914 21786
rect 6094 21734 6096 21786
rect 5850 21732 5856 21734
rect 5912 21732 5936 21734
rect 5992 21732 6016 21734
rect 6072 21732 6096 21734
rect 6152 21732 6158 21734
rect 5850 21723 6158 21732
rect 6380 21690 6408 22578
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6104 21010 6132 21286
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 5816 20936 5868 20942
rect 5736 20896 5816 20924
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5184 19502 5304 19530
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 388 18760 440 18766
rect 388 18702 440 18708
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 400 18465 428 18702
rect 2850 18524 3158 18533
rect 2850 18522 2856 18524
rect 2912 18522 2936 18524
rect 2992 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3158 18524
rect 2912 18470 2914 18522
rect 3094 18470 3096 18522
rect 2850 18468 2856 18470
rect 2912 18468 2936 18470
rect 2992 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3158 18470
rect 386 18456 442 18465
rect 2850 18459 3158 18468
rect 3620 18426 3648 18702
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 386 18391 442 18400
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3804 18358 3832 18566
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 4172 18086 4200 19110
rect 4350 19068 4658 19077
rect 4350 19066 4356 19068
rect 4412 19066 4436 19068
rect 4492 19066 4516 19068
rect 4572 19066 4596 19068
rect 4652 19066 4658 19068
rect 4412 19014 4414 19066
rect 4594 19014 4596 19066
rect 4350 19012 4356 19014
rect 4412 19012 4436 19014
rect 4492 19012 4516 19014
rect 4572 19012 4596 19014
rect 4652 19012 4658 19014
rect 4350 19003 4658 19012
rect 4724 18698 4752 19110
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 5092 18358 5120 18702
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 5184 18222 5212 19502
rect 5632 19440 5684 19446
rect 5632 19382 5684 19388
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5276 18834 5304 19246
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5276 18154 5304 18770
rect 5460 18426 5488 19110
rect 5644 18970 5672 19382
rect 5736 18986 5764 20896
rect 5816 20878 5868 20884
rect 5850 20700 6158 20709
rect 5850 20698 5856 20700
rect 5912 20698 5936 20700
rect 5992 20698 6016 20700
rect 6072 20698 6096 20700
rect 6152 20698 6158 20700
rect 5912 20646 5914 20698
rect 6094 20646 6096 20698
rect 5850 20644 5856 20646
rect 5912 20644 5936 20646
rect 5992 20644 6016 20646
rect 6072 20644 6096 20646
rect 6152 20644 6158 20646
rect 5850 20635 6158 20644
rect 5850 19612 6158 19621
rect 5850 19610 5856 19612
rect 5912 19610 5936 19612
rect 5992 19610 6016 19612
rect 6072 19610 6096 19612
rect 6152 19610 6158 19612
rect 5912 19558 5914 19610
rect 6094 19558 6096 19610
rect 5850 19556 5856 19558
rect 5912 19556 5936 19558
rect 5992 19556 6016 19558
rect 6072 19556 6096 19558
rect 6152 19556 6158 19558
rect 5850 19547 6158 19556
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5736 18958 5856 18986
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 1350 17980 1658 17989
rect 1350 17978 1356 17980
rect 1412 17978 1436 17980
rect 1492 17978 1516 17980
rect 1572 17978 1596 17980
rect 1652 17978 1658 17980
rect 1412 17926 1414 17978
rect 1594 17926 1596 17978
rect 1350 17924 1356 17926
rect 1412 17924 1436 17926
rect 1492 17924 1516 17926
rect 1572 17924 1596 17926
rect 1652 17924 1658 17926
rect 1350 17915 1658 17924
rect 4172 17678 4200 18022
rect 4350 17980 4658 17989
rect 4350 17978 4356 17980
rect 4412 17978 4436 17980
rect 4492 17978 4516 17980
rect 4572 17978 4596 17980
rect 4652 17978 4658 17980
rect 4412 17926 4414 17978
rect 4594 17926 4596 17978
rect 4350 17924 4356 17926
rect 4412 17924 4436 17926
rect 4492 17924 4516 17926
rect 4572 17924 4596 17926
rect 4652 17924 4658 17926
rect 4350 17915 4658 17924
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 5644 17610 5672 18022
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 2850 17436 3158 17445
rect 2850 17434 2856 17436
rect 2912 17434 2936 17436
rect 2992 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3158 17436
rect 2912 17382 2914 17434
rect 3094 17382 3096 17434
rect 2850 17380 2856 17382
rect 2912 17380 2936 17382
rect 2992 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3158 17382
rect 2850 17371 3158 17380
rect 5736 17338 5764 18958
rect 5828 18766 5856 18958
rect 6104 18834 6132 19246
rect 6288 18834 6316 20946
rect 6472 20398 6500 23462
rect 6564 23254 6592 23530
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6656 23066 6684 23122
rect 6564 23038 6684 23066
rect 6564 21078 6592 23038
rect 6644 22976 6696 22982
rect 6748 22930 6776 23666
rect 7024 23186 7052 24006
rect 7116 23866 7144 24142
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 6696 22924 6776 22930
rect 6644 22918 6776 22924
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6656 22902 6776 22918
rect 6748 22778 6776 22902
rect 6840 22778 6868 22918
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22094 6868 22510
rect 6656 22066 6868 22094
rect 6656 21486 6684 22066
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6748 21554 6776 21898
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6656 20924 6684 21422
rect 6564 20896 6684 20924
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 6472 19242 6500 20334
rect 6564 19310 6592 20896
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 19854 6684 20742
rect 6748 20466 6776 21490
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7024 21010 7052 21422
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7024 20602 7052 20946
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7116 20466 7144 20742
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7208 20058 7236 24754
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7350 24508 7658 24517
rect 7350 24506 7356 24508
rect 7412 24506 7436 24508
rect 7492 24506 7516 24508
rect 7572 24506 7596 24508
rect 7652 24506 7658 24508
rect 7412 24454 7414 24506
rect 7594 24454 7596 24506
rect 7350 24452 7356 24454
rect 7412 24452 7436 24454
rect 7492 24452 7516 24454
rect 7572 24452 7596 24454
rect 7652 24452 7658 24454
rect 7350 24443 7658 24452
rect 7288 24064 7340 24070
rect 7288 24006 7340 24012
rect 7300 23798 7328 24006
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7350 23420 7658 23429
rect 7350 23418 7356 23420
rect 7412 23418 7436 23420
rect 7492 23418 7516 23420
rect 7572 23418 7596 23420
rect 7652 23418 7658 23420
rect 7412 23366 7414 23418
rect 7594 23366 7596 23418
rect 7350 23364 7356 23366
rect 7412 23364 7436 23366
rect 7492 23364 7516 23366
rect 7572 23364 7596 23366
rect 7652 23364 7658 23366
rect 7350 23355 7658 23364
rect 7852 23254 7880 24686
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7944 23662 7972 24074
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7944 22574 7972 23598
rect 8312 23322 8340 23734
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8404 22710 8432 24006
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7350 22332 7658 22341
rect 7350 22330 7356 22332
rect 7412 22330 7436 22332
rect 7492 22330 7516 22332
rect 7572 22330 7596 22332
rect 7652 22330 7658 22332
rect 7412 22278 7414 22330
rect 7594 22278 7596 22330
rect 7350 22276 7356 22278
rect 7412 22276 7436 22278
rect 7492 22276 7516 22278
rect 7572 22276 7596 22278
rect 7652 22276 7658 22278
rect 7350 22267 7658 22276
rect 7944 22098 7972 22510
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 7748 22024 7800 22030
rect 7654 21992 7710 22001
rect 7748 21966 7800 21972
rect 7654 21927 7656 21936
rect 7708 21927 7710 21936
rect 7656 21898 7708 21904
rect 7350 21244 7658 21253
rect 7350 21242 7356 21244
rect 7412 21242 7436 21244
rect 7492 21242 7516 21244
rect 7572 21242 7596 21244
rect 7652 21242 7658 21244
rect 7412 21190 7414 21242
rect 7594 21190 7596 21242
rect 7350 21188 7356 21190
rect 7412 21188 7436 21190
rect 7492 21188 7516 21190
rect 7572 21188 7596 21190
rect 7652 21188 7658 21190
rect 7350 21179 7658 21188
rect 7760 20602 7788 21966
rect 7944 21486 7972 22034
rect 8024 21888 8076 21894
rect 8024 21830 8076 21836
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7944 20942 7972 21422
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 8036 20874 8064 21830
rect 8024 20868 8076 20874
rect 8024 20810 8076 20816
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 8588 20534 8616 20742
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 7350 20156 7658 20165
rect 7350 20154 7356 20156
rect 7412 20154 7436 20156
rect 7492 20154 7516 20156
rect 7572 20154 7596 20156
rect 7652 20154 7658 20156
rect 7412 20102 7414 20154
rect 7594 20102 7596 20154
rect 7350 20100 7356 20102
rect 7412 20100 7436 20102
rect 7492 20100 7516 20102
rect 7572 20100 7596 20102
rect 7652 20100 7658 20102
rect 7350 20091 7658 20100
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5850 18524 6158 18533
rect 5850 18522 5856 18524
rect 5912 18522 5936 18524
rect 5992 18522 6016 18524
rect 6072 18522 6096 18524
rect 6152 18522 6158 18524
rect 5912 18470 5914 18522
rect 6094 18470 6096 18522
rect 5850 18468 5856 18470
rect 5912 18468 5936 18470
rect 5992 18468 6016 18470
rect 6072 18468 6096 18470
rect 6152 18468 6158 18470
rect 5850 18459 6158 18468
rect 6380 18290 6408 19110
rect 6472 18290 6500 19178
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 5850 17436 6158 17445
rect 5850 17434 5856 17436
rect 5912 17434 5936 17436
rect 5992 17434 6016 17436
rect 6072 17434 6096 17436
rect 6152 17434 6158 17436
rect 5912 17382 5914 17434
rect 6094 17382 6096 17434
rect 5850 17380 5856 17382
rect 5912 17380 5936 17382
rect 5992 17380 6016 17382
rect 6072 17380 6096 17382
rect 6152 17380 6158 17382
rect 5850 17371 6158 17380
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 1350 16892 1658 16901
rect 1350 16890 1356 16892
rect 1412 16890 1436 16892
rect 1492 16890 1516 16892
rect 1572 16890 1596 16892
rect 1652 16890 1658 16892
rect 1412 16838 1414 16890
rect 1594 16838 1596 16890
rect 1350 16836 1356 16838
rect 1412 16836 1436 16838
rect 1492 16836 1516 16838
rect 1572 16836 1596 16838
rect 1652 16836 1658 16838
rect 1350 16827 1658 16836
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 1308 16448 1360 16454
rect 1306 16416 1308 16425
rect 1360 16416 1362 16425
rect 1306 16351 1362 16360
rect 2516 16250 2544 16458
rect 2792 16250 2820 16526
rect 2850 16348 3158 16357
rect 2850 16346 2856 16348
rect 2912 16346 2936 16348
rect 2992 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3158 16348
rect 2912 16294 2914 16346
rect 3094 16294 3096 16346
rect 2850 16292 2856 16294
rect 2912 16292 2936 16294
rect 2992 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3158 16294
rect 2850 16283 3158 16292
rect 3896 16250 3924 16594
rect 4264 16454 4292 17002
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4350 16892 4658 16901
rect 4350 16890 4356 16892
rect 4412 16890 4436 16892
rect 4492 16890 4516 16892
rect 4572 16890 4596 16892
rect 4652 16890 4658 16892
rect 4412 16838 4414 16890
rect 4594 16838 4596 16890
rect 4350 16836 4356 16838
rect 4412 16836 4436 16838
rect 4492 16836 4516 16838
rect 4572 16836 4596 16838
rect 4652 16836 4658 16838
rect 4350 16827 4658 16836
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 756 16108 808 16114
rect 756 16050 808 16056
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 768 15745 796 16050
rect 1350 15804 1658 15813
rect 1350 15802 1356 15804
rect 1412 15802 1436 15804
rect 1492 15802 1516 15804
rect 1572 15802 1596 15804
rect 1652 15802 1658 15804
rect 1412 15750 1414 15802
rect 1594 15750 1596 15802
rect 1350 15748 1356 15750
rect 1412 15748 1436 15750
rect 1492 15748 1516 15750
rect 1572 15748 1596 15750
rect 1652 15748 1658 15750
rect 754 15736 810 15745
rect 1350 15739 1658 15748
rect 754 15671 810 15680
rect 2240 15638 2268 16050
rect 2228 15632 2280 15638
rect 2228 15574 2280 15580
rect 2792 15570 2820 16186
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2884 15706 2912 16118
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 1216 15020 1268 15026
rect 1398 14991 1454 15000
rect 1216 14962 1268 14968
rect 754 14376 810 14385
rect 754 14311 810 14320
rect 768 14278 796 14311
rect 756 14272 808 14278
rect 756 14214 808 14220
rect 1228 13705 1256 14962
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 1350 14716 1658 14725
rect 1350 14714 1356 14716
rect 1412 14714 1436 14716
rect 1492 14714 1516 14716
rect 1572 14714 1596 14716
rect 1652 14714 1658 14716
rect 1412 14662 1414 14714
rect 1594 14662 1596 14714
rect 1350 14660 1356 14662
rect 1412 14660 1436 14662
rect 1492 14660 1516 14662
rect 1572 14660 1596 14662
rect 1652 14660 1658 14662
rect 1350 14651 1658 14660
rect 2700 14482 2728 14758
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1872 13938 1900 14214
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1214 13696 1270 13705
rect 1214 13631 1270 13640
rect 1350 13628 1658 13637
rect 1350 13626 1356 13628
rect 1412 13626 1436 13628
rect 1492 13626 1516 13628
rect 1572 13626 1596 13628
rect 1652 13626 1658 13628
rect 1412 13574 1414 13626
rect 1594 13574 1596 13626
rect 1350 13572 1356 13574
rect 1412 13572 1436 13574
rect 1492 13572 1516 13574
rect 1572 13572 1596 13574
rect 1652 13572 1658 13574
rect 1350 13563 1658 13572
rect 1688 13530 1716 13874
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 1306 13016 1362 13025
rect 1872 12986 1900 13194
rect 2608 12986 2636 13194
rect 1306 12951 1308 12960
rect 1360 12951 1362 12960
rect 1860 12980 1912 12986
rect 1308 12922 1360 12928
rect 1860 12922 1912 12928
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2700 12918 2728 14418
rect 2792 14006 2820 15506
rect 3528 15502 3556 15914
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15570 4200 15846
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 2850 15260 3158 15269
rect 2850 15258 2856 15260
rect 2912 15258 2936 15260
rect 2992 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3158 15260
rect 2912 15206 2914 15258
rect 3094 15206 3096 15258
rect 2850 15204 2856 15206
rect 2912 15204 2936 15206
rect 2992 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3158 15206
rect 2850 15195 3158 15204
rect 4172 15162 4200 15302
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 15094 4292 16390
rect 4448 16250 4476 16390
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4350 15804 4658 15813
rect 4350 15802 4356 15804
rect 4412 15802 4436 15804
rect 4492 15802 4516 15804
rect 4572 15802 4596 15804
rect 4652 15802 4658 15804
rect 4412 15750 4414 15802
rect 4594 15750 4596 15802
rect 4350 15748 4356 15750
rect 4412 15748 4436 15750
rect 4492 15748 4516 15750
rect 4572 15748 4596 15750
rect 4652 15748 4658 15750
rect 4350 15739 4658 15748
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4448 15026 4476 15506
rect 4724 15366 4752 15982
rect 4816 15502 4844 15982
rect 5092 15502 5120 16934
rect 5276 16590 5304 17274
rect 6564 17270 6592 19246
rect 6656 18358 6684 19314
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 5276 15162 5304 16118
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5460 15026 5488 16934
rect 5552 15910 5580 17138
rect 5644 16114 5672 17138
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5736 16658 5764 17002
rect 6472 16658 6500 17070
rect 6564 17066 6592 17206
rect 6748 17066 6776 18770
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6932 18222 6960 18702
rect 7024 18358 7052 19314
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18970 7144 19246
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7208 18426 7236 19110
rect 7350 19068 7658 19077
rect 7350 19066 7356 19068
rect 7412 19066 7436 19068
rect 7492 19066 7516 19068
rect 7572 19066 7596 19068
rect 7652 19066 7658 19068
rect 7412 19014 7414 19066
rect 7594 19014 7596 19066
rect 7350 19012 7356 19014
rect 7412 19012 7436 19014
rect 7492 19012 7516 19014
rect 7572 19012 7596 19014
rect 7652 19012 7658 19014
rect 7350 19003 7658 19012
rect 8680 18698 8708 24550
rect 8772 24206 8800 26982
rect 8956 26874 8984 26982
rect 9034 26924 9090 27324
rect 9678 26924 9734 27324
rect 10322 26924 10378 27324
rect 10966 26924 11022 27324
rect 11610 26924 11666 27324
rect 12254 26924 12310 27324
rect 12898 26924 12954 27324
rect 13542 26924 13598 27324
rect 14186 26924 14242 27324
rect 14830 26924 14886 27324
rect 15474 26924 15530 27324
rect 16118 26924 16174 27324
rect 18694 26924 18750 27324
rect 19338 26924 19394 27324
rect 19982 26924 20038 27324
rect 9048 26874 9076 26924
rect 8956 26846 9076 26874
rect 8850 25052 9158 25061
rect 8850 25050 8856 25052
rect 8912 25050 8936 25052
rect 8992 25050 9016 25052
rect 9072 25050 9096 25052
rect 9152 25050 9158 25052
rect 8912 24998 8914 25050
rect 9094 24998 9096 25050
rect 8850 24996 8856 24998
rect 8912 24996 8936 24998
rect 8992 24996 9016 24998
rect 9072 24996 9096 24998
rect 9152 24996 9158 24998
rect 8850 24987 9158 24996
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 9324 24614 9352 24822
rect 9692 24818 9720 26924
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9404 24608 9456 24614
rect 9404 24550 9456 24556
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8772 22030 8800 24006
rect 8850 23964 9158 23973
rect 8850 23962 8856 23964
rect 8912 23962 8936 23964
rect 8992 23962 9016 23964
rect 9072 23962 9096 23964
rect 9152 23962 9158 23964
rect 8912 23910 8914 23962
rect 9094 23910 9096 23962
rect 8850 23908 8856 23910
rect 8912 23908 8936 23910
rect 8992 23908 9016 23910
rect 9072 23908 9096 23910
rect 9152 23908 9158 23910
rect 8850 23899 9158 23908
rect 8850 22876 9158 22885
rect 8850 22874 8856 22876
rect 8912 22874 8936 22876
rect 8992 22874 9016 22876
rect 9072 22874 9096 22876
rect 9152 22874 9158 22876
rect 8912 22822 8914 22874
rect 9094 22822 9096 22874
rect 8850 22820 8856 22822
rect 8912 22820 8936 22822
rect 8992 22820 9016 22822
rect 9072 22820 9096 22822
rect 9152 22820 9158 22822
rect 8850 22811 9158 22820
rect 9232 22642 9260 24210
rect 9324 24206 9352 24550
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9324 22778 9352 24006
rect 9416 23186 9444 24550
rect 9508 23730 9536 24550
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9508 23066 9536 23122
rect 9416 23038 9536 23066
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9232 22166 9260 22578
rect 9416 22234 9444 23038
rect 9496 22976 9548 22982
rect 9600 22964 9628 24006
rect 9876 23866 9904 24074
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9968 23730 9996 24142
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 9548 22936 9628 22964
rect 9496 22918 9548 22924
rect 9508 22710 9536 22918
rect 9692 22778 9720 23666
rect 9968 22982 9996 23666
rect 10152 23526 10180 24686
rect 10336 24682 10364 26924
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10350 24508 10658 24517
rect 10350 24506 10356 24508
rect 10412 24506 10436 24508
rect 10492 24506 10516 24508
rect 10572 24506 10596 24508
rect 10652 24506 10658 24508
rect 10412 24454 10414 24506
rect 10594 24454 10596 24506
rect 10350 24452 10356 24454
rect 10412 24452 10436 24454
rect 10492 24452 10516 24454
rect 10572 24452 10596 24454
rect 10652 24452 10658 24454
rect 10350 24443 10658 24452
rect 10796 23730 10824 24686
rect 10980 24410 11008 26924
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23730 11376 24006
rect 11440 23866 11468 24686
rect 11520 24676 11572 24682
rect 11520 24618 11572 24624
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10350 23420 10658 23429
rect 10350 23418 10356 23420
rect 10412 23418 10436 23420
rect 10492 23418 10516 23420
rect 10572 23418 10596 23420
rect 10652 23418 10658 23420
rect 10412 23366 10414 23418
rect 10594 23366 10596 23418
rect 10350 23364 10356 23366
rect 10412 23364 10436 23366
rect 10492 23364 10516 23366
rect 10572 23364 10596 23366
rect 10652 23364 10658 23366
rect 10350 23355 10658 23364
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9496 22704 9548 22710
rect 9496 22646 9548 22652
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 9416 22094 9444 22170
rect 9416 22066 9536 22094
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 8850 21788 9158 21797
rect 8850 21786 8856 21788
rect 8912 21786 8936 21788
rect 8992 21786 9016 21788
rect 9072 21786 9096 21788
rect 9152 21786 9158 21788
rect 8912 21734 8914 21786
rect 9094 21734 9096 21786
rect 8850 21732 8856 21734
rect 8912 21732 8936 21734
rect 8992 21732 9016 21734
rect 9072 21732 9096 21734
rect 9152 21732 9158 21734
rect 8850 21723 9158 21732
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8864 21146 8892 21490
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 9232 20942 9260 21830
rect 9416 21622 9444 21966
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 8772 20058 8800 20878
rect 8850 20700 9158 20709
rect 8850 20698 8856 20700
rect 8912 20698 8936 20700
rect 8992 20698 9016 20700
rect 9072 20698 9096 20700
rect 9152 20698 9158 20700
rect 8912 20646 8914 20698
rect 9094 20646 9096 20698
rect 8850 20644 8856 20646
rect 8912 20644 8936 20646
rect 8992 20644 9016 20646
rect 9072 20644 9096 20646
rect 9152 20644 9158 20646
rect 8850 20635 9158 20644
rect 9324 20602 9352 20946
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8850 19612 9158 19621
rect 8850 19610 8856 19612
rect 8912 19610 8936 19612
rect 8992 19610 9016 19612
rect 9072 19610 9096 19612
rect 9152 19610 9158 19612
rect 8912 19558 8914 19610
rect 9094 19558 9096 19610
rect 8850 19556 8856 19558
rect 8912 19556 8936 19558
rect 8992 19556 9016 19558
rect 9072 19556 9096 19558
rect 9152 19556 9158 19558
rect 8850 19547 9158 19556
rect 9324 19310 9352 20538
rect 9416 19854 9444 21558
rect 9508 19922 9536 22066
rect 9968 21554 9996 22918
rect 10060 22642 10088 23122
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10350 22332 10658 22341
rect 10350 22330 10356 22332
rect 10412 22330 10436 22332
rect 10492 22330 10516 22332
rect 10572 22330 10596 22332
rect 10652 22330 10658 22332
rect 10412 22278 10414 22330
rect 10594 22278 10596 22330
rect 10350 22276 10356 22278
rect 10412 22276 10436 22278
rect 10492 22276 10516 22278
rect 10572 22276 10596 22278
rect 10652 22276 10658 22278
rect 10350 22267 10658 22276
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 9956 21548 10008 21554
rect 9876 21508 9956 21536
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9692 20618 9720 21422
rect 9600 20590 9720 20618
rect 9600 20534 9628 20590
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9876 20466 9904 21508
rect 9956 21490 10008 21496
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 21146 10180 21286
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10244 21026 10272 21830
rect 10336 21350 10364 21966
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10350 21244 10658 21253
rect 10350 21242 10356 21244
rect 10412 21242 10436 21244
rect 10492 21242 10516 21244
rect 10572 21242 10596 21244
rect 10652 21242 10658 21244
rect 10412 21190 10414 21242
rect 10594 21190 10596 21242
rect 10350 21188 10356 21190
rect 10412 21188 10436 21190
rect 10492 21188 10516 21190
rect 10572 21188 10596 21190
rect 10652 21188 10658 21190
rect 10350 21179 10658 21188
rect 10244 20998 10364 21026
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9692 20058 9720 20402
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9416 19514 9444 19654
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9508 18766 9536 19858
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9692 18834 9720 19314
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6932 17882 6960 18158
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7116 17678 7144 18022
rect 7350 17980 7658 17989
rect 7350 17978 7356 17980
rect 7412 17978 7436 17980
rect 7492 17978 7516 17980
rect 7572 17978 7596 17980
rect 7652 17978 7658 17980
rect 7412 17926 7414 17978
rect 7594 17926 7596 17978
rect 7350 17924 7356 17926
rect 7412 17924 7436 17926
rect 7492 17924 7516 17926
rect 7572 17924 7596 17926
rect 7652 17924 7658 17926
rect 7350 17915 7658 17924
rect 7760 17882 7788 18634
rect 8680 18358 8708 18634
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 8772 18426 8800 18566
rect 8850 18524 9158 18533
rect 8850 18522 8856 18524
rect 8912 18522 8936 18524
rect 8992 18522 9016 18524
rect 9072 18522 9096 18524
rect 9152 18522 9158 18524
rect 8912 18470 8914 18522
rect 9094 18470 9096 18522
rect 8850 18468 8856 18470
rect 8912 18468 8936 18470
rect 8992 18468 9016 18470
rect 9072 18468 9096 18470
rect 9152 18468 9158 18470
rect 8850 18459 9158 18468
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6748 16810 6776 17002
rect 6656 16782 6776 16810
rect 6840 16794 6868 17274
rect 6828 16788 6880 16794
rect 6656 16726 6684 16782
rect 6828 16730 6880 16736
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 7208 16658 7236 17614
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7760 17338 7788 17546
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 7350 16892 7658 16901
rect 7350 16890 7356 16892
rect 7412 16890 7436 16892
rect 7492 16890 7516 16892
rect 7572 16890 7596 16892
rect 7652 16890 7658 16892
rect 7412 16838 7414 16890
rect 7594 16838 7596 16890
rect 7350 16836 7356 16838
rect 7412 16836 7436 16838
rect 7492 16836 7516 16838
rect 7572 16836 7596 16838
rect 7652 16836 7658 16838
rect 7350 16827 7658 16836
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 5850 16348 6158 16357
rect 5850 16346 5856 16348
rect 5912 16346 5936 16348
rect 5992 16346 6016 16348
rect 6072 16346 6096 16348
rect 6152 16346 6158 16348
rect 5912 16294 5914 16346
rect 6094 16294 6096 16346
rect 5850 16292 5856 16294
rect 5912 16292 5936 16294
rect 5992 16292 6016 16294
rect 6072 16292 6096 16294
rect 6152 16292 6158 16294
rect 5850 16283 6158 16292
rect 6288 16182 6316 16526
rect 6472 16250 6500 16594
rect 8036 16590 8064 16934
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 6288 15706 6316 16118
rect 8312 16114 8340 18226
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8404 17134 8432 18022
rect 8680 17542 8708 18294
rect 9324 18290 9352 18566
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8680 17338 8708 17478
rect 8850 17436 9158 17445
rect 8850 17434 8856 17436
rect 8912 17434 8936 17436
rect 8992 17434 9016 17436
rect 9072 17434 9096 17436
rect 9152 17434 9158 17436
rect 8912 17382 8914 17434
rect 9094 17382 9096 17434
rect 8850 17380 8856 17382
rect 8912 17380 8936 17382
rect 8992 17380 9016 17382
rect 9072 17380 9096 17382
rect 9152 17380 9158 17382
rect 8850 17371 9158 17380
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 9508 17134 9536 18702
rect 9600 17746 9628 18702
rect 9692 18290 9720 18770
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9692 17270 9720 18226
rect 9968 17954 9996 20878
rect 10336 20534 10364 20998
rect 10324 20528 10376 20534
rect 10324 20470 10376 20476
rect 10350 20156 10658 20165
rect 10350 20154 10356 20156
rect 10412 20154 10436 20156
rect 10492 20154 10516 20156
rect 10572 20154 10596 20156
rect 10652 20154 10658 20156
rect 10412 20102 10414 20154
rect 10594 20102 10596 20154
rect 10350 20100 10356 20102
rect 10412 20100 10436 20102
rect 10492 20100 10516 20102
rect 10572 20100 10596 20102
rect 10652 20100 10658 20102
rect 10350 20091 10658 20100
rect 10704 19310 10732 23054
rect 10796 19922 10824 23666
rect 11242 23624 11298 23633
rect 11242 23559 11298 23568
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10888 23118 10916 23462
rect 11256 23254 11284 23559
rect 11440 23254 11468 23802
rect 11532 23610 11560 24618
rect 11624 24614 11652 26924
rect 11850 25052 12158 25061
rect 11850 25050 11856 25052
rect 11912 25050 11936 25052
rect 11992 25050 12016 25052
rect 12072 25050 12096 25052
rect 12152 25050 12158 25052
rect 11912 24998 11914 25050
rect 12094 24998 12096 25050
rect 11850 24996 11856 24998
rect 11912 24996 11936 24998
rect 11992 24996 12016 24998
rect 12072 24996 12096 24998
rect 12152 24996 12158 24998
rect 11850 24987 12158 24996
rect 12268 24750 12296 26924
rect 12912 24818 12940 26924
rect 13556 24818 13584 26924
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 12452 24410 12480 24754
rect 12900 24676 12952 24682
rect 12900 24618 12952 24624
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11532 23582 11652 23610
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 11532 22778 11560 23462
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11520 22024 11572 22030
rect 11242 21992 11298 22001
rect 11520 21966 11572 21972
rect 11242 21927 11298 21936
rect 10876 21004 10928 21010
rect 10876 20946 10928 20952
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10888 19802 10916 20946
rect 11256 20942 11284 21927
rect 11532 21690 11560 21966
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11348 21010 11376 21286
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11244 20936 11296 20942
rect 11072 20896 11244 20924
rect 11072 20754 11100 20896
rect 11244 20878 11296 20884
rect 10796 19774 10916 19802
rect 10980 20726 11100 20754
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10244 18834 10272 19178
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10350 19068 10658 19077
rect 10350 19066 10356 19068
rect 10412 19066 10436 19068
rect 10492 19066 10516 19068
rect 10572 19066 10596 19068
rect 10652 19066 10658 19068
rect 10412 19014 10414 19066
rect 10594 19014 10596 19066
rect 10350 19012 10356 19014
rect 10412 19012 10436 19014
rect 10492 19012 10516 19014
rect 10572 19012 10596 19014
rect 10652 19012 10658 19014
rect 10350 19003 10658 19012
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10244 18358 10272 18770
rect 10704 18698 10732 19110
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10796 18578 10824 19774
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10704 18550 10824 18578
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 9784 17926 9996 17954
rect 10350 17980 10658 17989
rect 10350 17978 10356 17980
rect 10412 17978 10436 17980
rect 10492 17978 10516 17980
rect 10572 17978 10596 17980
rect 10652 17978 10658 17980
rect 10412 17926 10414 17978
rect 10594 17926 10596 17978
rect 9784 17678 9812 17926
rect 10350 17924 10356 17926
rect 10412 17924 10436 17926
rect 10492 17924 10516 17926
rect 10572 17924 10596 17926
rect 10652 17924 10658 17926
rect 10350 17915 10658 17924
rect 10704 17746 10732 18550
rect 10888 18426 10916 19246
rect 10980 18698 11008 20726
rect 11164 19922 11192 20742
rect 11256 20466 11284 20742
rect 11348 20466 11376 20946
rect 11440 20874 11468 21354
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11440 20602 11468 20810
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11256 19854 11284 20402
rect 11532 20346 11560 21422
rect 11440 20318 11560 20346
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10888 17746 10916 18362
rect 10980 18329 11008 18634
rect 10966 18320 11022 18329
rect 10966 18255 11022 18264
rect 11072 17882 11100 19314
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9864 17672 9916 17678
rect 10244 17626 10272 17682
rect 9864 17614 9916 17620
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9508 16726 9536 17070
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9692 16590 9720 17070
rect 9784 16794 9812 17614
rect 9876 17134 9904 17614
rect 10152 17598 10272 17626
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 10152 16998 10180 17598
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9600 16402 9628 16526
rect 9600 16374 9720 16402
rect 8850 16348 9158 16357
rect 8850 16346 8856 16348
rect 8912 16346 8936 16348
rect 8992 16346 9016 16348
rect 9072 16346 9096 16348
rect 9152 16346 9158 16348
rect 8912 16294 8914 16346
rect 9094 16294 9096 16346
rect 8850 16292 8856 16294
rect 8912 16292 8936 16294
rect 8992 16292 9016 16294
rect 9072 16292 9096 16294
rect 9152 16292 9158 16294
rect 8850 16283 9158 16292
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 5850 15260 6158 15269
rect 5850 15258 5856 15260
rect 5912 15258 5936 15260
rect 5992 15258 6016 15260
rect 6072 15258 6096 15260
rect 6152 15258 6158 15260
rect 5912 15206 5914 15258
rect 6094 15206 6096 15258
rect 5850 15204 5856 15206
rect 5912 15204 5936 15206
rect 5992 15204 6016 15206
rect 6072 15204 6096 15206
rect 6152 15204 6158 15206
rect 5850 15195 6158 15204
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 14414 2912 14758
rect 2976 14482 3004 14962
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2850 14172 3158 14181
rect 2850 14170 2856 14172
rect 2912 14170 2936 14172
rect 2992 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3158 14172
rect 2912 14118 2914 14170
rect 3094 14118 3096 14170
rect 2850 14116 2856 14118
rect 2912 14116 2936 14118
rect 2992 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3158 14118
rect 2850 14107 3158 14116
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2792 12918 2820 13942
rect 2850 13084 3158 13093
rect 2850 13082 2856 13084
rect 2912 13082 2936 13084
rect 2992 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3158 13084
rect 2912 13030 2914 13082
rect 3094 13030 3096 13082
rect 2850 13028 2856 13030
rect 2912 13028 2936 13030
rect 2992 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3158 13030
rect 2850 13019 3158 13028
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 1350 12540 1658 12549
rect 1350 12538 1356 12540
rect 1412 12538 1436 12540
rect 1492 12538 1516 12540
rect 1572 12538 1596 12540
rect 1652 12538 1658 12540
rect 1412 12486 1414 12538
rect 1594 12486 1596 12538
rect 1350 12484 1356 12486
rect 1412 12484 1436 12486
rect 1492 12484 1516 12486
rect 1572 12484 1596 12486
rect 1652 12484 1658 12486
rect 1350 12475 1658 12484
rect 386 12336 442 12345
rect 386 12271 442 12280
rect 400 12238 428 12271
rect 388 12232 440 12238
rect 388 12174 440 12180
rect 2850 11996 3158 12005
rect 2850 11994 2856 11996
rect 2912 11994 2936 11996
rect 2992 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3158 11996
rect 2912 11942 2914 11994
rect 3094 11942 3096 11994
rect 2850 11940 2856 11942
rect 2912 11940 2936 11942
rect 2992 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3158 11942
rect 2850 11931 3158 11940
rect 3344 11778 3372 14962
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3436 12238 3464 13942
rect 3528 13938 3556 14214
rect 4172 14074 4200 14214
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4080 13954 4108 14010
rect 4264 13954 4292 14894
rect 4350 14716 4658 14725
rect 4350 14714 4356 14716
rect 4412 14714 4436 14716
rect 4492 14714 4516 14716
rect 4572 14714 4596 14716
rect 4652 14714 4658 14716
rect 4412 14662 4414 14714
rect 4594 14662 4596 14714
rect 4350 14660 4356 14662
rect 4412 14660 4436 14662
rect 4492 14660 4516 14662
rect 4572 14660 4596 14662
rect 4652 14660 4658 14662
rect 4350 14651 4658 14660
rect 4908 14482 4936 14894
rect 6656 14890 6684 15982
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7350 15804 7658 15813
rect 7350 15802 7356 15804
rect 7412 15802 7436 15804
rect 7492 15802 7516 15804
rect 7572 15802 7596 15804
rect 7652 15802 7658 15804
rect 7412 15750 7414 15802
rect 7594 15750 7596 15802
rect 7350 15748 7356 15750
rect 7412 15748 7436 15750
rect 7492 15748 7516 15750
rect 7572 15748 7596 15750
rect 7652 15748 7658 15750
rect 7350 15739 7658 15748
rect 7944 15638 7972 15846
rect 9692 15706 9720 16374
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 3516 13932 3568 13938
rect 4080 13926 4292 13954
rect 3516 13874 3568 13880
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4172 13394 4200 13670
rect 4264 13530 4292 13926
rect 4632 13802 4660 14350
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4350 13628 4658 13637
rect 4350 13626 4356 13628
rect 4412 13626 4436 13628
rect 4492 13626 4516 13628
rect 4572 13626 4596 13628
rect 4652 13626 4658 13628
rect 4412 13574 4414 13626
rect 4594 13574 4596 13626
rect 4350 13572 4356 13574
rect 4412 13572 4436 13574
rect 4492 13572 4516 13574
rect 4572 13572 4596 13574
rect 4652 13572 4658 13574
rect 4350 13563 4658 13572
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3896 12986 3924 13262
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 4356 13138 4384 13330
rect 4724 13326 4752 13466
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4816 13138 4844 13738
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3988 12850 4016 13126
rect 4356 13110 4844 13138
rect 4356 12866 4384 13110
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4172 12838 4384 12866
rect 4528 12844 4580 12850
rect 3896 12753 3924 12786
rect 3882 12744 3938 12753
rect 3882 12679 3938 12688
rect 3988 12238 4016 12786
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 388 11756 440 11762
rect 388 11698 440 11704
rect 3240 11756 3292 11762
rect 3344 11750 3556 11778
rect 3240 11698 3292 11704
rect 400 11665 428 11698
rect 386 11656 442 11665
rect 386 11591 442 11600
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1350 11452 1658 11461
rect 1350 11450 1356 11452
rect 1412 11450 1436 11452
rect 1492 11450 1516 11452
rect 1572 11450 1596 11452
rect 1652 11450 1658 11452
rect 1412 11398 1414 11450
rect 1594 11398 1596 11450
rect 1350 11396 1356 11398
rect 1412 11396 1436 11398
rect 1492 11396 1516 11398
rect 1572 11396 1596 11398
rect 1652 11396 1658 11398
rect 1350 11387 1658 11396
rect 1688 11150 1716 11562
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 11150 2820 11494
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 3252 11082 3280 11698
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1860 11008 1912 11014
rect 1544 10976 1546 10985
rect 1860 10950 1912 10956
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 1490 10911 1546 10920
rect 1872 10577 1900 10950
rect 2148 10742 2176 10950
rect 2850 10908 3158 10917
rect 2850 10906 2856 10908
rect 2912 10906 2936 10908
rect 2992 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3158 10908
rect 2912 10854 2914 10906
rect 3094 10854 3096 10906
rect 2850 10852 2856 10854
rect 2912 10852 2936 10854
rect 2992 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3158 10854
rect 2850 10843 3158 10852
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 1858 10568 1914 10577
rect 1858 10503 1914 10512
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1350 10364 1658 10373
rect 1350 10362 1356 10364
rect 1412 10362 1436 10364
rect 1492 10362 1516 10364
rect 1572 10362 1596 10364
rect 1652 10362 1658 10364
rect 1412 10310 1414 10362
rect 1594 10310 1596 10362
rect 1350 10308 1356 10310
rect 1412 10308 1436 10310
rect 1492 10308 1516 10310
rect 1572 10308 1596 10310
rect 1652 10308 1658 10310
rect 1350 10299 1658 10308
rect 1872 9994 1900 10406
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1780 9722 1808 9930
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 386 9616 442 9625
rect 386 9551 388 9560
rect 440 9551 442 9560
rect 388 9522 440 9528
rect 1350 9276 1658 9285
rect 1350 9274 1356 9276
rect 1412 9274 1436 9276
rect 1492 9274 1516 9276
rect 1572 9274 1596 9276
rect 1652 9274 1658 9276
rect 1412 9222 1414 9274
rect 1594 9222 1596 9274
rect 1350 9220 1356 9222
rect 1412 9220 1436 9222
rect 1492 9220 1516 9222
rect 1572 9220 1596 9222
rect 1652 9220 1658 9222
rect 1350 9211 1658 9220
rect 388 8968 440 8974
rect 386 8936 388 8945
rect 440 8936 442 8945
rect 386 8871 442 8880
rect 1872 8430 1900 9930
rect 2850 9820 3158 9829
rect 2850 9818 2856 9820
rect 2912 9818 2936 9820
rect 2992 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3158 9820
rect 2912 9766 2914 9818
rect 3094 9766 3096 9818
rect 2850 9764 2856 9766
rect 2912 9764 2936 9766
rect 2992 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3158 9766
rect 2850 9755 3158 9764
rect 3252 9722 3280 11018
rect 3344 11014 3372 11630
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 11150 3464 11494
rect 3528 11218 3556 11750
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3620 11082 3648 11222
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10810 3372 10950
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 9722 3464 10610
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 10198 3556 10542
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8566 2268 8774
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1216 8356 1268 8362
rect 1216 8298 1268 8304
rect 1228 8265 1256 8298
rect 1214 8256 1270 8265
rect 1214 8191 1270 8200
rect 1350 8188 1658 8197
rect 1350 8186 1356 8188
rect 1412 8186 1436 8188
rect 1492 8186 1516 8188
rect 1572 8186 1596 8188
rect 1652 8186 1658 8188
rect 1412 8134 1414 8186
rect 1594 8134 1596 8186
rect 1350 8132 1356 8134
rect 1412 8132 1436 8134
rect 1492 8132 1516 8134
rect 1572 8132 1596 8134
rect 1652 8132 1658 8134
rect 1350 8123 1658 8132
rect 1872 7886 1900 8366
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 2792 7342 2820 9386
rect 3712 9110 3740 11154
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3804 10062 3832 11086
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3896 9926 3924 10542
rect 4068 10532 4120 10538
rect 4172 10520 4200 12838
rect 4528 12786 4580 12792
rect 4540 12730 4568 12786
rect 4264 12702 4568 12730
rect 4264 12442 4292 12702
rect 4350 12540 4658 12549
rect 4350 12538 4356 12540
rect 4412 12538 4436 12540
rect 4492 12538 4516 12540
rect 4572 12538 4596 12540
rect 4652 12538 4658 12540
rect 4412 12486 4414 12538
rect 4594 12486 4596 12538
rect 4350 12484 4356 12486
rect 4412 12484 4436 12486
rect 4492 12484 4516 12486
rect 4572 12484 4596 12486
rect 4652 12484 4658 12486
rect 4350 12475 4658 12484
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4908 11694 4936 14418
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5276 13734 5304 13806
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4350 11452 4658 11461
rect 4350 11450 4356 11452
rect 4412 11450 4436 11452
rect 4492 11450 4516 11452
rect 4572 11450 4596 11452
rect 4652 11450 4658 11452
rect 4412 11398 4414 11450
rect 4594 11398 4596 11450
rect 4350 11396 4356 11398
rect 4412 11396 4436 11398
rect 4492 11396 4516 11398
rect 4572 11396 4596 11398
rect 4652 11396 4658 11398
rect 4350 11387 4658 11396
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10674 4292 10950
rect 5000 10690 5028 13330
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5092 11014 5120 11630
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10810 5120 10950
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4908 10662 5028 10690
rect 4908 10606 4936 10662
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4120 10492 4200 10520
rect 4068 10474 4120 10480
rect 4172 10266 4200 10492
rect 4350 10364 4658 10373
rect 4350 10362 4356 10364
rect 4412 10362 4436 10364
rect 4492 10362 4516 10364
rect 4572 10362 4596 10364
rect 4652 10362 4658 10364
rect 4412 10310 4414 10362
rect 4594 10310 4596 10362
rect 4350 10308 4356 10310
rect 4412 10308 4436 10310
rect 4492 10308 4516 10310
rect 4572 10308 4596 10310
rect 4652 10308 4658 10310
rect 4350 10299 4658 10308
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9586 3924 9862
rect 4172 9654 4200 10066
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 4350 9276 4658 9285
rect 4350 9274 4356 9276
rect 4412 9274 4436 9276
rect 4492 9274 4516 9276
rect 4572 9274 4596 9276
rect 4652 9274 4658 9276
rect 4412 9222 4414 9274
rect 4594 9222 4596 9274
rect 4350 9220 4356 9222
rect 4412 9220 4436 9222
rect 4492 9220 4516 9222
rect 4572 9220 4596 9222
rect 4652 9220 4658 9222
rect 4350 9211 4658 9220
rect 4724 9160 4752 10542
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4816 9674 4844 10202
rect 4908 9994 4936 10406
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4816 9646 4936 9674
rect 4356 9132 4752 9160
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2850 8732 3158 8741
rect 2850 8730 2856 8732
rect 2912 8730 2936 8732
rect 2992 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3158 8732
rect 2912 8678 2914 8730
rect 3094 8678 3096 8730
rect 2850 8676 2856 8678
rect 2912 8676 2936 8678
rect 2992 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3158 8678
rect 2850 8667 3158 8676
rect 3252 8634 3280 8910
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7818 3372 8230
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 2850 7644 3158 7653
rect 2850 7642 2856 7644
rect 2912 7642 2936 7644
rect 2992 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3158 7644
rect 2912 7590 2914 7642
rect 3094 7590 3096 7642
rect 2850 7588 2856 7590
rect 2912 7588 2936 7590
rect 2992 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3158 7590
rect 2850 7579 3158 7588
rect 3528 7546 3556 8434
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3804 7886 3832 8026
rect 4172 7886 4200 8774
rect 4356 8498 4384 9132
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8498 4660 8910
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4908 8430 4936 9646
rect 5276 9518 5304 13670
rect 5368 12986 5396 13806
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5552 12646 5580 14214
rect 5736 13530 5764 14350
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 5850 14172 6158 14181
rect 5850 14170 5856 14172
rect 5912 14170 5936 14172
rect 5992 14170 6016 14172
rect 6072 14170 6096 14172
rect 6152 14170 6158 14172
rect 5912 14118 5914 14170
rect 6094 14118 6096 14170
rect 5850 14116 5856 14118
rect 5912 14116 5936 14118
rect 5992 14116 6016 14118
rect 6072 14116 6096 14118
rect 6152 14116 6158 14118
rect 5850 14107 6158 14116
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 6196 13326 6224 14214
rect 6564 14074 6592 14350
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6656 13734 6684 14826
rect 7024 14278 7052 15370
rect 7576 15162 7604 15370
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14414 7236 14758
rect 7350 14716 7658 14725
rect 7350 14714 7356 14716
rect 7412 14714 7436 14716
rect 7492 14714 7516 14716
rect 7572 14714 7596 14716
rect 7652 14714 7658 14716
rect 7412 14662 7414 14714
rect 7594 14662 7596 14714
rect 7350 14660 7356 14662
rect 7412 14660 7436 14662
rect 7492 14660 7516 14662
rect 7572 14660 7596 14662
rect 7652 14660 7658 14662
rect 7350 14651 7658 14660
rect 7760 14618 7788 15438
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6932 14074 6960 14214
rect 7024 14074 7052 14214
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 7024 13326 7052 14010
rect 7116 13734 7144 14350
rect 7392 13938 7420 14554
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7944 13870 7972 15574
rect 8128 15366 8156 15574
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13530 7144 13670
rect 7350 13628 7658 13637
rect 7350 13626 7356 13628
rect 7412 13626 7436 13628
rect 7492 13626 7516 13628
rect 7572 13626 7596 13628
rect 7652 13626 7658 13628
rect 7412 13574 7414 13626
rect 7594 13574 7596 13626
rect 7350 13572 7356 13574
rect 7412 13572 7436 13574
rect 7492 13572 7516 13574
rect 7572 13572 7596 13574
rect 7652 13572 7658 13574
rect 7350 13563 7658 13572
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7852 13326 7880 13738
rect 8128 13394 8156 15302
rect 8220 15162 8248 15302
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8312 14890 8340 15506
rect 9692 15502 9720 15642
rect 9968 15502 9996 15914
rect 10152 15638 10180 16934
rect 10244 16794 10272 17138
rect 10350 16892 10658 16901
rect 10350 16890 10356 16892
rect 10412 16890 10436 16892
rect 10492 16890 10516 16892
rect 10572 16890 10596 16892
rect 10652 16890 10658 16892
rect 10412 16838 10414 16890
rect 10594 16838 10596 16890
rect 10350 16836 10356 16838
rect 10412 16836 10436 16838
rect 10492 16836 10516 16838
rect 10572 16836 10596 16838
rect 10652 16836 10658 16838
rect 10350 16827 10658 16836
rect 10796 16794 10824 17274
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 11072 16658 11100 17478
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 15994 11008 16526
rect 10704 15966 11008 15994
rect 10350 15804 10658 15813
rect 10350 15802 10356 15804
rect 10412 15802 10436 15804
rect 10492 15802 10516 15804
rect 10572 15802 10596 15804
rect 10652 15802 10658 15804
rect 10412 15750 10414 15802
rect 10594 15750 10596 15802
rect 10350 15748 10356 15750
rect 10412 15748 10436 15750
rect 10492 15748 10516 15750
rect 10572 15748 10596 15750
rect 10652 15748 10658 15750
rect 10350 15739 10658 15748
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 8850 15260 9158 15269
rect 8850 15258 8856 15260
rect 8912 15258 8936 15260
rect 8992 15258 9016 15260
rect 9072 15258 9096 15260
rect 9152 15258 9158 15260
rect 8912 15206 8914 15258
rect 9094 15206 9096 15258
rect 8850 15204 8856 15206
rect 8912 15204 8936 15206
rect 8992 15204 9016 15206
rect 9072 15204 9096 15206
rect 9152 15204 9158 15206
rect 8850 15195 9158 15204
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 8312 14074 8340 14826
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14482 9168 14758
rect 9416 14618 9444 14962
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 5850 13084 6158 13093
rect 5850 13082 5856 13084
rect 5912 13082 5936 13084
rect 5992 13082 6016 13084
rect 6072 13082 6096 13084
rect 6152 13082 6158 13084
rect 5912 13030 5914 13082
rect 6094 13030 6096 13082
rect 5850 13028 5856 13030
rect 5912 13028 5936 13030
rect 5992 13028 6016 13030
rect 6072 13028 6096 13030
rect 6152 13028 6158 13030
rect 5850 13019 6158 13028
rect 6182 12744 6238 12753
rect 6182 12679 6238 12688
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5850 11996 6158 12005
rect 5850 11994 5856 11996
rect 5912 11994 5936 11996
rect 5992 11994 6016 11996
rect 6072 11994 6096 11996
rect 6152 11994 6158 11996
rect 5912 11942 5914 11994
rect 6094 11942 6096 11994
rect 5850 11940 5856 11942
rect 5912 11940 5936 11942
rect 5992 11940 6016 11942
rect 6072 11940 6096 11942
rect 6152 11940 6158 11942
rect 5850 11931 6158 11940
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5368 10606 5396 11086
rect 5460 10810 5488 11698
rect 5850 10908 6158 10917
rect 5850 10906 5856 10908
rect 5912 10906 5936 10908
rect 5992 10906 6016 10908
rect 6072 10906 6096 10908
rect 6152 10906 6158 10908
rect 5912 10854 5914 10906
rect 6094 10854 6096 10906
rect 5850 10852 5856 10854
rect 5912 10852 5936 10854
rect 5992 10852 6016 10854
rect 6072 10852 6096 10854
rect 6152 10852 6158 10854
rect 5850 10843 6158 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 6196 10742 6224 12679
rect 6656 12646 6684 13262
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7392 12986 7420 13126
rect 7852 12986 7880 13126
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 8404 12850 8432 13806
rect 8588 13258 8616 13806
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8680 12714 8708 13262
rect 8772 12918 8800 14350
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8850 14172 9158 14181
rect 8850 14170 8856 14172
rect 8912 14170 8936 14172
rect 8992 14170 9016 14172
rect 9072 14170 9096 14172
rect 9152 14170 9158 14172
rect 8912 14118 8914 14170
rect 9094 14118 9096 14170
rect 8850 14116 8856 14118
rect 8912 14116 8936 14118
rect 8992 14116 9016 14118
rect 9072 14116 9096 14118
rect 9152 14116 9158 14118
rect 8850 14107 9158 14116
rect 9232 14074 9260 14282
rect 9508 14074 9536 15098
rect 9600 14482 9628 15302
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10060 14618 10088 14962
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 10244 14414 10272 15302
rect 10350 14716 10658 14725
rect 10350 14714 10356 14716
rect 10412 14714 10436 14716
rect 10492 14714 10516 14716
rect 10572 14714 10596 14716
rect 10652 14714 10658 14716
rect 10412 14662 10414 14714
rect 10594 14662 10596 14714
rect 10350 14660 10356 14662
rect 10412 14660 10436 14662
rect 10492 14660 10516 14662
rect 10572 14660 10596 14662
rect 10652 14660 10658 14662
rect 10350 14651 10658 14660
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 8850 13084 9158 13093
rect 8850 13082 8856 13084
rect 8912 13082 8936 13084
rect 8992 13082 9016 13084
rect 9072 13082 9096 13084
rect 9152 13082 9158 13084
rect 8912 13030 8914 13082
rect 9094 13030 9096 13082
rect 8850 13028 8856 13030
rect 8912 13028 8936 13030
rect 8992 13028 9016 13030
rect 9072 13028 9096 13030
rect 9152 13028 9158 13030
rect 8850 13019 9158 13028
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6184 10736 6236 10742
rect 6182 10704 6184 10713
rect 6236 10704 6238 10713
rect 6182 10639 6238 10648
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5368 10062 5396 10542
rect 5644 10266 5672 10542
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5276 9042 5304 9454
rect 5552 9110 5580 9454
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5644 9042 5672 10202
rect 5850 9820 6158 9829
rect 5850 9818 5856 9820
rect 5912 9818 5936 9820
rect 5992 9818 6016 9820
rect 6072 9818 6096 9820
rect 6152 9818 6158 9820
rect 5912 9766 5914 9818
rect 6094 9766 6096 9818
rect 5850 9764 5856 9766
rect 5912 9764 5936 9766
rect 5992 9764 6016 9766
rect 6072 9764 6096 9766
rect 6152 9764 6158 9766
rect 5850 9755 6158 9764
rect 6380 9722 6408 10610
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9178 5856 9522
rect 6472 9178 6500 11018
rect 6656 9654 6684 12582
rect 7350 12540 7658 12549
rect 7350 12538 7356 12540
rect 7412 12538 7436 12540
rect 7492 12538 7516 12540
rect 7572 12538 7596 12540
rect 7652 12538 7658 12540
rect 7412 12486 7414 12538
rect 7594 12486 7596 12538
rect 7350 12484 7356 12486
rect 7412 12484 7436 12486
rect 7492 12484 7516 12486
rect 7572 12484 7596 12486
rect 7652 12484 7658 12486
rect 7350 12475 7658 12484
rect 8680 12434 8708 12650
rect 8588 12406 8708 12434
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 10062 6776 10406
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6840 9654 6868 11494
rect 7350 11452 7658 11461
rect 7350 11450 7356 11452
rect 7412 11450 7436 11452
rect 7492 11450 7516 11452
rect 7572 11450 7596 11452
rect 7652 11450 7658 11452
rect 7412 11398 7414 11450
rect 7594 11398 7596 11450
rect 7350 11396 7356 11398
rect 7412 11396 7436 11398
rect 7492 11396 7516 11398
rect 7572 11396 7596 11398
rect 7652 11396 7658 11398
rect 7350 11387 7658 11396
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10810 7052 11018
rect 7760 11014 7788 11630
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11354 8156 11494
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7760 10674 7788 10950
rect 8220 10713 8248 11018
rect 8206 10704 8262 10713
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7748 10668 7800 10674
rect 8206 10639 8262 10648
rect 7748 10610 7800 10616
rect 7668 10554 7696 10610
rect 7208 10538 7788 10554
rect 7196 10532 7788 10538
rect 7248 10526 7788 10532
rect 7196 10474 7248 10480
rect 7350 10364 7658 10373
rect 7350 10362 7356 10364
rect 7412 10362 7436 10364
rect 7492 10362 7516 10364
rect 7572 10362 7596 10364
rect 7652 10362 7658 10364
rect 7412 10310 7414 10362
rect 7594 10310 7596 10362
rect 7350 10308 7356 10310
rect 7412 10308 7436 10310
rect 7492 10308 7516 10310
rect 7572 10308 7596 10310
rect 7652 10308 7658 10310
rect 7350 10299 7658 10308
rect 7760 10266 7788 10526
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9722 7144 9998
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 8220 9654 8248 10639
rect 8312 10470 8340 11698
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8496 11014 8524 11630
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10674 8524 10950
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8588 10606 8616 12406
rect 8772 12238 8800 12854
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12238 9444 12582
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8680 11354 8708 12174
rect 8850 11996 9158 12005
rect 8850 11994 8856 11996
rect 8912 11994 8936 11996
rect 8992 11994 9016 11996
rect 9072 11994 9096 11996
rect 9152 11994 9158 11996
rect 8912 11942 8914 11994
rect 9094 11942 9096 11994
rect 8850 11940 8856 11942
rect 8912 11940 8936 11942
rect 8992 11940 9016 11942
rect 9072 11940 9096 11942
rect 9152 11940 9158 11942
rect 8850 11931 9158 11940
rect 9232 11830 9260 12174
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9416 11762 9444 12038
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8942 11112 8998 11121
rect 8942 11047 8944 11056
rect 8996 11047 8998 11056
rect 8944 11018 8996 11024
rect 8850 10908 9158 10917
rect 8850 10906 8856 10908
rect 8912 10906 8936 10908
rect 8992 10906 9016 10908
rect 9072 10906 9096 10908
rect 9152 10906 9158 10908
rect 8912 10854 8914 10906
rect 9094 10854 9096 10906
rect 8850 10852 8856 10854
rect 8912 10852 8936 10854
rect 8992 10852 9016 10854
rect 9072 10852 9096 10854
rect 9152 10852 9158 10854
rect 8850 10843 9158 10852
rect 9416 10810 9444 11494
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9508 10690 9536 14010
rect 10704 13938 10732 15966
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10980 15570 11008 15846
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11060 14816 11112 14822
rect 11164 14804 11192 18226
rect 11440 17746 11468 20318
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 19990 11560 20198
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11624 19514 11652 23582
rect 11716 20058 11744 24074
rect 11850 23964 12158 23973
rect 11850 23962 11856 23964
rect 11912 23962 11936 23964
rect 11992 23962 12016 23964
rect 12072 23962 12096 23964
rect 12152 23962 12158 23964
rect 11912 23910 11914 23962
rect 12094 23910 12096 23962
rect 11850 23908 11856 23910
rect 11912 23908 11936 23910
rect 11992 23908 12016 23910
rect 12072 23908 12096 23910
rect 12152 23908 12158 23910
rect 11850 23899 12158 23908
rect 12268 23746 12296 24142
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 12176 23718 12296 23746
rect 11900 23186 11928 23666
rect 12176 23322 12204 23718
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 12268 23118 12296 23598
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12440 23112 12492 23118
rect 12544 23100 12572 24006
rect 12728 23798 12756 24006
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12492 23072 12572 23100
rect 12440 23054 12492 23060
rect 11850 22876 12158 22885
rect 11850 22874 11856 22876
rect 11912 22874 11936 22876
rect 11992 22874 12016 22876
rect 12072 22874 12096 22876
rect 12152 22874 12158 22876
rect 11912 22822 11914 22874
rect 12094 22822 12096 22874
rect 11850 22820 11856 22822
rect 11912 22820 11936 22822
rect 11992 22820 12016 22822
rect 12072 22820 12096 22822
rect 12152 22820 12158 22822
rect 11850 22811 12158 22820
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 11850 21788 12158 21797
rect 11850 21786 11856 21788
rect 11912 21786 11936 21788
rect 11992 21786 12016 21788
rect 12072 21786 12096 21788
rect 12152 21786 12158 21788
rect 11912 21734 11914 21786
rect 12094 21734 12096 21786
rect 11850 21732 11856 21734
rect 11912 21732 11936 21734
rect 11992 21732 12016 21734
rect 12072 21732 12096 21734
rect 12152 21732 12158 21734
rect 11850 21723 12158 21732
rect 12544 20942 12572 21830
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 11850 20700 12158 20709
rect 11850 20698 11856 20700
rect 11912 20698 11936 20700
rect 11992 20698 12016 20700
rect 12072 20698 12096 20700
rect 12152 20698 12158 20700
rect 11912 20646 11914 20698
rect 12094 20646 12096 20698
rect 11850 20644 11856 20646
rect 11912 20644 11936 20646
rect 11992 20644 12016 20646
rect 12072 20644 12096 20646
rect 12152 20644 12158 20646
rect 11850 20635 12158 20644
rect 12728 20534 12756 21830
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11850 19612 12158 19621
rect 11850 19610 11856 19612
rect 11912 19610 11936 19612
rect 11992 19610 12016 19612
rect 12072 19610 12096 19612
rect 12152 19610 12158 19612
rect 11912 19558 11914 19610
rect 12094 19558 12096 19610
rect 11850 19556 11856 19558
rect 11912 19556 11936 19558
rect 11992 19556 12016 19558
rect 12072 19556 12096 19558
rect 12152 19556 12158 19558
rect 11850 19547 12158 19556
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11716 18222 11744 18702
rect 11850 18524 12158 18533
rect 11850 18522 11856 18524
rect 11912 18522 11936 18524
rect 11992 18522 12016 18524
rect 12072 18522 12096 18524
rect 12152 18522 12158 18524
rect 11912 18470 11914 18522
rect 12094 18470 12096 18522
rect 11850 18468 11856 18470
rect 11912 18468 11936 18470
rect 11992 18468 12016 18470
rect 12072 18468 12096 18470
rect 12152 18468 12158 18470
rect 11850 18459 12158 18468
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 12360 18170 12388 19178
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18358 12572 18566
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12728 18290 12756 19110
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 11716 17746 11744 18158
rect 12360 18142 12480 18170
rect 12452 18086 12480 18142
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11348 17338 11376 17614
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11440 16794 11468 17682
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 17338 11560 17478
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11716 17270 11744 17682
rect 11992 17678 12020 18022
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 12452 17490 12480 18022
rect 12268 17462 12480 17490
rect 11850 17436 12158 17445
rect 11850 17434 11856 17436
rect 11912 17434 11936 17436
rect 11992 17434 12016 17436
rect 12072 17434 12096 17436
rect 12152 17434 12158 17436
rect 11912 17382 11914 17434
rect 12094 17382 12096 17434
rect 11850 17380 11856 17382
rect 11912 17380 11936 17382
rect 11992 17380 12016 17382
rect 12072 17380 12096 17382
rect 12152 17380 12158 17382
rect 11850 17371 12158 17380
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 12268 17202 12296 17462
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11850 16348 12158 16357
rect 11850 16346 11856 16348
rect 11912 16346 11936 16348
rect 11992 16346 12016 16348
rect 12072 16346 12096 16348
rect 12152 16346 12158 16348
rect 11912 16294 11914 16346
rect 12094 16294 12096 16346
rect 11850 16292 11856 16294
rect 11912 16292 11936 16294
rect 11992 16292 12016 16294
rect 12072 16292 12096 16294
rect 12152 16292 12158 16294
rect 11850 16283 12158 16292
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11256 15162 11284 15982
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11256 14958 11284 15098
rect 11348 15026 11376 15302
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11112 14776 11192 14804
rect 11060 14758 11112 14764
rect 11072 14278 11100 14758
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10350 13628 10658 13637
rect 10350 13626 10356 13628
rect 10412 13626 10436 13628
rect 10492 13626 10516 13628
rect 10572 13626 10596 13628
rect 10652 13626 10658 13628
rect 10412 13574 10414 13626
rect 10594 13574 10596 13626
rect 10350 13572 10356 13574
rect 10412 13572 10436 13574
rect 10492 13572 10516 13574
rect 10572 13572 10596 13574
rect 10652 13572 10658 13574
rect 10350 13563 10658 13572
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 12442 10180 12718
rect 10350 12540 10658 12549
rect 10350 12538 10356 12540
rect 10412 12538 10436 12540
rect 10492 12538 10516 12540
rect 10572 12538 10596 12540
rect 10652 12538 10658 12540
rect 10412 12486 10414 12538
rect 10594 12486 10596 12538
rect 10350 12484 10356 12486
rect 10412 12484 10436 12486
rect 10492 12484 10516 12486
rect 10572 12484 10596 12486
rect 10652 12484 10658 12486
rect 10350 12475 10658 12484
rect 10140 12436 10192 12442
rect 10704 12434 10732 13874
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10704 12406 10824 12434
rect 10140 12378 10192 12384
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9600 11082 9628 11766
rect 10152 11762 10180 12378
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10796 11778 10824 12406
rect 10888 11898 10916 13262
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11072 12306 11100 12718
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11164 11898 11192 13262
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12918 11376 13126
rect 11440 12986 11468 15506
rect 11532 15094 11560 15574
rect 11716 15502 11744 15846
rect 11900 15570 11928 16050
rect 12360 15570 12388 17206
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12728 16522 12756 17138
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 11850 15260 12158 15269
rect 11850 15258 11856 15260
rect 11912 15258 11936 15260
rect 11992 15258 12016 15260
rect 12072 15258 12096 15260
rect 12152 15258 12158 15260
rect 11912 15206 11914 15258
rect 12094 15206 12096 15258
rect 11850 15204 11856 15206
rect 11912 15204 11936 15206
rect 11992 15204 12016 15206
rect 12072 15204 12096 15206
rect 12152 15204 12158 15206
rect 11850 15195 12158 15204
rect 12452 15162 12480 15370
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 12728 15026 12756 16458
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14346 11560 14758
rect 11808 14550 11836 14962
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11850 14172 12158 14181
rect 11850 14170 11856 14172
rect 11912 14170 11936 14172
rect 11992 14170 12016 14172
rect 12072 14170 12096 14172
rect 12152 14170 12158 14172
rect 11912 14118 11914 14170
rect 12094 14118 12096 14170
rect 11850 14116 11856 14118
rect 11912 14116 11936 14118
rect 11992 14116 12016 14118
rect 12072 14116 12096 14118
rect 12152 14116 12158 14118
rect 11850 14107 12158 14116
rect 12452 13530 12480 14486
rect 12532 14000 12584 14006
rect 12530 13968 12532 13977
rect 12584 13968 12586 13977
rect 12530 13903 12586 13912
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11428 12980 11480 12986
rect 11480 12940 11560 12968
rect 11428 12922 11480 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11440 12442 11468 12786
rect 11532 12646 11560 12940
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10152 11150 10180 11698
rect 10350 11452 10658 11461
rect 10350 11450 10356 11452
rect 10412 11450 10436 11452
rect 10492 11450 10516 11452
rect 10572 11450 10596 11452
rect 10652 11450 10658 11452
rect 10412 11398 10414 11450
rect 10594 11398 10596 11450
rect 10350 11396 10356 11398
rect 10412 11396 10436 11398
rect 10492 11396 10516 11398
rect 10572 11396 10596 11398
rect 10652 11396 10658 11398
rect 10350 11387 10658 11396
rect 10704 11218 10732 11766
rect 10796 11750 11192 11778
rect 11164 11694 11192 11750
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11072 11354 11100 11630
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9416 10662 9536 10690
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 10266 8708 10406
rect 8772 10266 8800 10542
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 6656 9466 6684 9590
rect 6828 9512 6880 9518
rect 6656 9460 6828 9466
rect 6656 9454 6880 9460
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 6656 9438 6868 9454
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 6656 8974 6684 9318
rect 7350 9276 7658 9285
rect 7350 9274 7356 9276
rect 7412 9274 7436 9276
rect 7492 9274 7516 9276
rect 7572 9274 7596 9276
rect 7652 9274 7658 9276
rect 7412 9222 7414 9274
rect 7594 9222 7596 9274
rect 7350 9220 7356 9222
rect 7412 9220 7436 9222
rect 7492 9220 7516 9222
rect 7572 9220 7596 9222
rect 7652 9220 7658 9222
rect 7350 9211 7658 9220
rect 7944 9042 7972 9454
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 8312 8838 8340 9930
rect 8404 9586 8432 9930
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8680 8974 8708 10202
rect 8850 9820 9158 9829
rect 8850 9818 8856 9820
rect 8912 9818 8936 9820
rect 8992 9818 9016 9820
rect 9072 9818 9096 9820
rect 9152 9818 9158 9820
rect 8912 9766 8914 9818
rect 9094 9766 9096 9818
rect 8850 9764 8856 9766
rect 8912 9764 8936 9766
rect 8992 9764 9016 9766
rect 9072 9764 9096 9766
rect 9152 9764 9158 9766
rect 8850 9755 9158 9764
rect 9324 9722 9352 10610
rect 9416 10606 9444 10662
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9220 9648 9272 9654
rect 9416 9602 9444 10542
rect 9600 10130 9628 11018
rect 11256 10674 11284 12174
rect 11440 11626 11468 12174
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11440 11218 11468 11562
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 10350 10364 10658 10373
rect 10350 10362 10356 10364
rect 10412 10362 10436 10364
rect 10492 10362 10516 10364
rect 10572 10362 10596 10364
rect 10652 10362 10658 10364
rect 10412 10310 10414 10362
rect 10594 10310 10596 10362
rect 10350 10308 10356 10310
rect 10412 10308 10436 10310
rect 10492 10308 10516 10310
rect 10572 10308 10596 10310
rect 10652 10308 10658 10310
rect 10350 10299 10658 10308
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10520 9722 10548 9930
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 9220 9590 9272 9596
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 4528 8424 4580 8430
rect 4896 8424 4948 8430
rect 4580 8372 4752 8378
rect 4528 8366 4752 8372
rect 4896 8366 4948 8372
rect 4540 8350 4752 8366
rect 4350 8188 4658 8197
rect 4350 8186 4356 8188
rect 4412 8186 4436 8188
rect 4492 8186 4516 8188
rect 4572 8186 4596 8188
rect 4652 8186 4658 8188
rect 4412 8134 4414 8186
rect 4594 8134 4596 8186
rect 4350 8132 4356 8134
rect 4412 8132 4436 8134
rect 4492 8132 4516 8134
rect 4572 8132 4596 8134
rect 4652 8132 4658 8134
rect 4350 8123 4658 8132
rect 4344 8016 4396 8022
rect 4264 7964 4344 7970
rect 4724 7970 4752 8350
rect 4908 8294 4936 8366
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4396 7964 4752 7970
rect 4264 7942 4752 7964
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3988 7478 4016 7686
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 1350 7100 1658 7109
rect 1350 7098 1356 7100
rect 1412 7098 1436 7100
rect 1492 7098 1516 7100
rect 1572 7098 1596 7100
rect 1652 7098 1658 7100
rect 1412 7046 1414 7098
rect 1594 7046 1596 7098
rect 1350 7044 1356 7046
rect 1412 7044 1436 7046
rect 1492 7044 1516 7046
rect 1572 7044 1596 7046
rect 1652 7044 1658 7046
rect 1350 7035 1658 7044
rect 2884 7002 2912 7278
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 4264 6866 4292 7942
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7206 4384 7822
rect 5000 7818 5028 8774
rect 5850 8732 6158 8741
rect 5850 8730 5856 8732
rect 5912 8730 5936 8732
rect 5992 8730 6016 8732
rect 6072 8730 6096 8732
rect 6152 8730 6158 8732
rect 5912 8678 5914 8730
rect 6094 8678 6096 8730
rect 5850 8676 5856 8678
rect 5912 8676 5936 8678
rect 5992 8676 6016 8678
rect 6072 8676 6096 8678
rect 6152 8676 6158 8678
rect 5850 8667 6158 8676
rect 6380 8634 6408 8774
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5552 7886 5580 8366
rect 5736 8022 5764 8366
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5540 7880 5592 7886
rect 6932 7834 6960 8230
rect 7350 8188 7658 8197
rect 7350 8186 7356 8188
rect 7412 8186 7436 8188
rect 7492 8186 7516 8188
rect 7572 8186 7596 8188
rect 7652 8186 7658 8188
rect 7412 8134 7414 8186
rect 7594 8134 7596 8186
rect 7350 8132 7356 8134
rect 7412 8132 7436 8134
rect 7492 8132 7516 8134
rect 7572 8132 7596 8134
rect 7652 8132 7658 8134
rect 7350 8123 7658 8132
rect 8036 8090 8064 8434
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7886 7972 7958
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7932 7880 7984 7886
rect 5540 7822 5592 7828
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5000 7410 5028 7754
rect 5552 7546 5580 7822
rect 6840 7806 6960 7834
rect 7852 7828 7932 7834
rect 7852 7822 7984 7828
rect 7748 7812 7800 7818
rect 5850 7644 6158 7653
rect 5850 7642 5856 7644
rect 5912 7642 5936 7644
rect 5992 7642 6016 7644
rect 6072 7642 6096 7644
rect 6152 7642 6158 7644
rect 5912 7590 5914 7642
rect 6094 7590 6096 7642
rect 5850 7588 5856 7590
rect 5912 7588 5936 7590
rect 5992 7588 6016 7590
rect 6072 7588 6096 7590
rect 6152 7588 6158 7590
rect 5850 7579 6158 7588
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 6840 7342 6868 7806
rect 7748 7754 7800 7760
rect 7852 7806 7972 7822
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4350 7100 4658 7109
rect 4350 7098 4356 7100
rect 4412 7098 4436 7100
rect 4492 7098 4516 7100
rect 4572 7098 4596 7100
rect 4652 7098 4658 7100
rect 4412 7046 4414 7098
rect 4594 7046 4596 7098
rect 4350 7044 4356 7046
rect 4412 7044 4436 7046
rect 4492 7044 4516 7046
rect 4572 7044 4596 7046
rect 4652 7044 4658 7046
rect 4350 7035 4658 7044
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 2850 6556 3158 6565
rect 2850 6554 2856 6556
rect 2912 6554 2936 6556
rect 2992 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3158 6556
rect 2912 6502 2914 6554
rect 3094 6502 3096 6554
rect 2850 6500 2856 6502
rect 2912 6500 2936 6502
rect 2992 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3158 6502
rect 2850 6491 3158 6500
rect 1350 6012 1658 6021
rect 1350 6010 1356 6012
rect 1412 6010 1436 6012
rect 1492 6010 1516 6012
rect 1572 6010 1596 6012
rect 1652 6010 1658 6012
rect 1412 5958 1414 6010
rect 1594 5958 1596 6010
rect 1350 5956 1356 5958
rect 1412 5956 1436 5958
rect 1492 5956 1516 5958
rect 1572 5956 1596 5958
rect 1652 5956 1658 5958
rect 1350 5947 1658 5956
rect 4350 6012 4658 6021
rect 4350 6010 4356 6012
rect 4412 6010 4436 6012
rect 4492 6010 4516 6012
rect 4572 6010 4596 6012
rect 4652 6010 4658 6012
rect 4412 5958 4414 6010
rect 4594 5958 4596 6010
rect 4350 5956 4356 5958
rect 4412 5956 4436 5958
rect 4492 5956 4516 5958
rect 4572 5956 4596 5958
rect 4652 5956 4658 5958
rect 4350 5947 4658 5956
rect 4724 5710 4752 7142
rect 6196 6798 6224 7278
rect 6932 6866 6960 7686
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5850 6556 6158 6565
rect 5850 6554 5856 6556
rect 5912 6554 5936 6556
rect 5992 6554 6016 6556
rect 6072 6554 6096 6556
rect 6152 6554 6158 6556
rect 5912 6502 5914 6554
rect 6094 6502 6096 6554
rect 5850 6500 5856 6502
rect 5912 6500 5936 6502
rect 5992 6500 6016 6502
rect 6072 6500 6096 6502
rect 6152 6500 6158 6502
rect 5850 6491 6158 6500
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 2850 5468 3158 5477
rect 2850 5466 2856 5468
rect 2912 5466 2936 5468
rect 2992 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3158 5468
rect 2912 5414 2914 5466
rect 3094 5414 3096 5466
rect 2850 5412 2856 5414
rect 2912 5412 2936 5414
rect 2992 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3158 5414
rect 2850 5403 3158 5412
rect 1350 4924 1658 4933
rect 1350 4922 1356 4924
rect 1412 4922 1436 4924
rect 1492 4922 1516 4924
rect 1572 4922 1596 4924
rect 1652 4922 1658 4924
rect 1412 4870 1414 4922
rect 1594 4870 1596 4922
rect 1350 4868 1356 4870
rect 1412 4868 1436 4870
rect 1492 4868 1516 4870
rect 1572 4868 1596 4870
rect 1652 4868 1658 4870
rect 1350 4859 1658 4868
rect 4350 4924 4658 4933
rect 4350 4922 4356 4924
rect 4412 4922 4436 4924
rect 4492 4922 4516 4924
rect 4572 4922 4596 4924
rect 4652 4922 4658 4924
rect 4412 4870 4414 4922
rect 4594 4870 4596 4922
rect 4350 4868 4356 4870
rect 4412 4868 4436 4870
rect 4492 4868 4516 4870
rect 4572 4868 4596 4870
rect 4652 4868 4658 4870
rect 4350 4859 4658 4868
rect 2850 4380 3158 4389
rect 2850 4378 2856 4380
rect 2912 4378 2936 4380
rect 2992 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3158 4380
rect 2912 4326 2914 4378
rect 3094 4326 3096 4378
rect 2850 4324 2856 4326
rect 2912 4324 2936 4326
rect 2992 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3158 4326
rect 2850 4315 3158 4324
rect 1350 3836 1658 3845
rect 1350 3834 1356 3836
rect 1412 3834 1436 3836
rect 1492 3834 1516 3836
rect 1572 3834 1596 3836
rect 1652 3834 1658 3836
rect 1412 3782 1414 3834
rect 1594 3782 1596 3834
rect 1350 3780 1356 3782
rect 1412 3780 1436 3782
rect 1492 3780 1516 3782
rect 1572 3780 1596 3782
rect 1652 3780 1658 3782
rect 1350 3771 1658 3780
rect 4350 3836 4658 3845
rect 4350 3834 4356 3836
rect 4412 3834 4436 3836
rect 4492 3834 4516 3836
rect 4572 3834 4596 3836
rect 4652 3834 4658 3836
rect 4412 3782 4414 3834
rect 4594 3782 4596 3834
rect 4350 3780 4356 3782
rect 4412 3780 4436 3782
rect 4492 3780 4516 3782
rect 4572 3780 4596 3782
rect 4652 3780 4658 3782
rect 4350 3771 4658 3780
rect 4724 3602 4752 5646
rect 5644 5370 5672 5714
rect 5850 5468 6158 5477
rect 5850 5466 5856 5468
rect 5912 5466 5936 5468
rect 5992 5466 6016 5468
rect 6072 5466 6096 5468
rect 6152 5466 6158 5468
rect 5912 5414 5914 5466
rect 6094 5414 6096 5466
rect 5850 5412 5856 5414
rect 5912 5412 5936 5414
rect 5992 5412 6016 5414
rect 6072 5412 6096 5414
rect 6152 5412 6158 5414
rect 5850 5403 6158 5412
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4690 5856 5102
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4146 5764 4422
rect 5850 4380 6158 4389
rect 5850 4378 5856 4380
rect 5912 4378 5936 4380
rect 5992 4378 6016 4380
rect 6072 4378 6096 4380
rect 6152 4378 6158 4380
rect 5912 4326 5914 4378
rect 6094 4326 6096 4378
rect 5850 4324 5856 4326
rect 5912 4324 5936 4326
rect 5992 4324 6016 4326
rect 6072 4324 6096 4326
rect 6152 4324 6158 4326
rect 5850 4315 6158 4324
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3602 5580 3878
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 2850 3292 3158 3301
rect 2850 3290 2856 3292
rect 2912 3290 2936 3292
rect 2992 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3158 3292
rect 2912 3238 2914 3290
rect 3094 3238 3096 3290
rect 2850 3236 2856 3238
rect 2912 3236 2936 3238
rect 2992 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3158 3238
rect 2850 3227 3158 3236
rect 5850 3292 6158 3301
rect 5850 3290 5856 3292
rect 5912 3290 5936 3292
rect 5992 3290 6016 3292
rect 6072 3290 6096 3292
rect 6152 3290 6158 3292
rect 5912 3238 5914 3290
rect 6094 3238 6096 3290
rect 5850 3236 5856 3238
rect 5912 3236 5936 3238
rect 5992 3236 6016 3238
rect 6072 3236 6096 3238
rect 6152 3236 6158 3238
rect 5850 3227 6158 3236
rect 6196 3058 6224 6734
rect 7208 6730 7236 7414
rect 7350 7100 7658 7109
rect 7350 7098 7356 7100
rect 7412 7098 7436 7100
rect 7492 7098 7516 7100
rect 7572 7098 7596 7100
rect 7652 7098 7658 7100
rect 7412 7046 7414 7098
rect 7594 7046 7596 7098
rect 7350 7044 7356 7046
rect 7412 7044 7436 7046
rect 7492 7044 7516 7046
rect 7572 7044 7596 7046
rect 7652 7044 7658 7046
rect 7350 7035 7658 7044
rect 7760 7002 7788 7754
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7852 6934 7880 7806
rect 7840 6928 7892 6934
rect 7760 6876 7840 6882
rect 7760 6870 7892 6876
rect 7760 6854 7880 6870
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 5642 7236 6666
rect 7350 6012 7658 6021
rect 7350 6010 7356 6012
rect 7412 6010 7436 6012
rect 7492 6010 7516 6012
rect 7572 6010 7596 6012
rect 7652 6010 7658 6012
rect 7412 5958 7414 6010
rect 7594 5958 7596 6010
rect 7350 5956 7356 5958
rect 7412 5956 7436 5958
rect 7492 5956 7516 5958
rect 7572 5956 7596 5958
rect 7652 5956 7658 5958
rect 7350 5947 7658 5956
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 6748 5302 6776 5578
rect 6840 5370 6868 5578
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6288 4146 6316 4422
rect 6656 4146 6684 5170
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 1350 2748 1658 2757
rect 1350 2746 1356 2748
rect 1412 2746 1436 2748
rect 1492 2746 1516 2748
rect 1572 2746 1596 2748
rect 1652 2746 1658 2748
rect 1412 2694 1414 2746
rect 1594 2694 1596 2746
rect 1350 2692 1356 2694
rect 1412 2692 1436 2694
rect 1492 2692 1516 2694
rect 1572 2692 1596 2694
rect 1652 2692 1658 2694
rect 1350 2683 1658 2692
rect 4350 2748 4658 2757
rect 4350 2746 4356 2748
rect 4412 2746 4436 2748
rect 4492 2746 4516 2748
rect 4572 2746 4596 2748
rect 4652 2746 4658 2748
rect 4412 2694 4414 2746
rect 4594 2694 4596 2746
rect 4350 2692 4356 2694
rect 4412 2692 4436 2694
rect 4492 2692 4516 2694
rect 4572 2692 4596 2694
rect 4652 2692 4658 2694
rect 4350 2683 4658 2692
rect 6748 2446 6776 5238
rect 7024 5234 7052 5510
rect 7392 5302 7420 5646
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7760 5234 7788 6854
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6338 8064 6598
rect 8128 6458 8156 7890
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8220 7546 8248 7754
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7342 8340 8774
rect 8850 8732 9158 8741
rect 8850 8730 8856 8732
rect 8912 8730 8936 8732
rect 8992 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9158 8732
rect 8912 8678 8914 8730
rect 9094 8678 9096 8730
rect 8850 8676 8856 8678
rect 8912 8676 8936 8678
rect 8992 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9158 8678
rect 8850 8667 9158 8676
rect 9232 8498 9260 9590
rect 9324 9574 9444 9602
rect 10140 9580 10192 9586
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 8864 7954 8892 8434
rect 9232 8090 9260 8434
rect 9324 8430 9352 9574
rect 10140 9522 10192 9528
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 8850 7644 9158 7653
rect 8850 7642 8856 7644
rect 8912 7642 8936 7644
rect 8992 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9158 7644
rect 8912 7590 8914 7642
rect 9094 7590 9096 7642
rect 8850 7588 8856 7590
rect 8912 7588 8936 7590
rect 8992 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9158 7590
rect 8850 7579 9158 7588
rect 9232 7410 9260 7822
rect 9324 7750 9352 8366
rect 9416 8294 9444 8978
rect 9508 8906 9536 9454
rect 9692 9178 9720 9454
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9508 7886 9536 8842
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8484 7404 8536 7410
rect 8852 7404 8904 7410
rect 8484 7346 8536 7352
rect 8772 7364 8852 7392
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8404 6662 8432 7346
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8036 6310 8156 6338
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 6840 4622 6868 5102
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4690 7236 5034
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7350 4924 7658 4933
rect 7350 4922 7356 4924
rect 7412 4922 7436 4924
rect 7492 4922 7516 4924
rect 7572 4922 7596 4924
rect 7652 4922 7658 4924
rect 7412 4870 7414 4922
rect 7594 4870 7596 4922
rect 7350 4868 7356 4870
rect 7412 4868 7436 4870
rect 7492 4868 7516 4870
rect 7572 4868 7596 4870
rect 7652 4868 7658 4870
rect 7350 4859 7658 4868
rect 7760 4758 7788 4966
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7852 4690 7880 5102
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6840 4282 6868 4558
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6932 4078 6960 4626
rect 7944 4554 7972 5238
rect 8036 5030 8064 5578
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7300 4282 7328 4422
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6840 3602 6868 4014
rect 7350 3836 7658 3845
rect 7350 3834 7356 3836
rect 7412 3834 7436 3836
rect 7492 3834 7516 3836
rect 7572 3834 7596 3836
rect 7652 3834 7658 3836
rect 7412 3782 7414 3834
rect 7594 3782 7596 3834
rect 7350 3780 7356 3782
rect 7412 3780 7436 3782
rect 7492 3780 7516 3782
rect 7572 3780 7596 3782
rect 7652 3780 7658 3782
rect 7350 3771 7658 3780
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 7760 3534 7788 4422
rect 7944 4146 7972 4490
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8036 3754 8064 4966
rect 7944 3726 8064 3754
rect 7944 3670 7972 3726
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7300 2938 7328 3402
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 3194 7604 3334
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7944 3126 7972 3606
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7208 2910 7328 2938
rect 7208 2650 7236 2910
rect 7300 2854 7328 2910
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7350 2748 7658 2757
rect 7350 2746 7356 2748
rect 7412 2746 7436 2748
rect 7492 2746 7516 2748
rect 7572 2746 7596 2748
rect 7652 2746 7658 2748
rect 7412 2694 7414 2746
rect 7594 2694 7596 2746
rect 7350 2692 7356 2694
rect 7412 2692 7436 2694
rect 7492 2692 7516 2694
rect 7572 2692 7596 2694
rect 7652 2692 7658 2694
rect 7350 2683 7658 2692
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 8036 2582 8064 3606
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8128 2446 8156 6310
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 5302 8432 6190
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8220 4826 8248 5102
rect 8496 5098 8524 7346
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 6730 8616 7142
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8588 5234 8616 6666
rect 8680 5370 8708 6802
rect 8772 5370 8800 7364
rect 8852 7346 8904 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 7002 9168 7142
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9232 6730 9260 7346
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 8850 6556 9158 6565
rect 8850 6554 8856 6556
rect 8912 6554 8936 6556
rect 8992 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9158 6556
rect 8912 6502 8914 6554
rect 9094 6502 9096 6554
rect 8850 6500 8856 6502
rect 8912 6500 8936 6502
rect 8992 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9158 6502
rect 8850 6491 9158 6500
rect 9324 6322 9352 7346
rect 9508 7342 9536 7822
rect 9600 7410 9628 8978
rect 10152 8634 10180 9522
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10350 9276 10658 9285
rect 10350 9274 10356 9276
rect 10412 9274 10436 9276
rect 10492 9274 10516 9276
rect 10572 9274 10596 9276
rect 10652 9274 10658 9276
rect 10412 9222 10414 9274
rect 10594 9222 10596 9274
rect 10350 9220 10356 9222
rect 10412 9220 10436 9222
rect 10492 9220 10516 9222
rect 10572 9220 10596 9222
rect 10652 9220 10658 9222
rect 10350 9211 10658 9220
rect 10796 9042 10824 9318
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6322 9536 7278
rect 10060 6798 10088 8502
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 8022 10180 8230
rect 10350 8188 10658 8197
rect 10350 8186 10356 8188
rect 10412 8186 10436 8188
rect 10492 8186 10516 8188
rect 10572 8186 10596 8188
rect 10652 8186 10658 8188
rect 10412 8134 10414 8186
rect 10594 8134 10596 8186
rect 10350 8132 10356 8134
rect 10412 8132 10436 8134
rect 10492 8132 10516 8134
rect 10572 8132 10596 8134
rect 10652 8132 10658 8134
rect 10350 8123 10658 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10350 7100 10658 7109
rect 10350 7098 10356 7100
rect 10412 7098 10436 7100
rect 10492 7098 10516 7100
rect 10572 7098 10596 7100
rect 10652 7098 10658 7100
rect 10412 7046 10414 7098
rect 10594 7046 10596 7098
rect 10350 7044 10356 7046
rect 10412 7044 10436 7046
rect 10492 7044 10516 7046
rect 10572 7044 10596 7046
rect 10652 7044 10658 7046
rect 10350 7035 10658 7044
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9140 5710 9168 6258
rect 9692 6118 9720 6598
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5710 9720 6054
rect 9784 5914 9812 6666
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9876 5914 9904 6190
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10060 5710 10088 6598
rect 11072 6458 11100 9930
rect 11532 9178 11560 12378
rect 11716 11898 11744 13126
rect 11850 13084 12158 13093
rect 11850 13082 11856 13084
rect 11912 13082 11936 13084
rect 11992 13082 12016 13084
rect 12072 13082 12096 13084
rect 12152 13082 12158 13084
rect 11912 13030 11914 13082
rect 12094 13030 12096 13082
rect 11850 13028 11856 13030
rect 11912 13028 11936 13030
rect 11992 13028 12016 13030
rect 12072 13028 12096 13030
rect 12152 13028 12158 13030
rect 11850 13019 12158 13028
rect 12360 12986 12388 13262
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11808 12374 11836 12650
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 12360 12306 12388 12922
rect 12728 12434 12756 14962
rect 12820 14414 12848 15846
rect 12912 15366 12940 24618
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 13096 22778 13124 24074
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13188 21690 13216 21966
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13280 19514 13308 24550
rect 13350 24508 13658 24517
rect 13350 24506 13356 24508
rect 13412 24506 13436 24508
rect 13492 24506 13516 24508
rect 13572 24506 13596 24508
rect 13652 24506 13658 24508
rect 13412 24454 13414 24506
rect 13594 24454 13596 24506
rect 13350 24452 13356 24454
rect 13412 24452 13436 24454
rect 13492 24452 13516 24454
rect 13572 24452 13596 24454
rect 13652 24452 13658 24454
rect 13350 24443 13658 24452
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13350 23420 13658 23429
rect 13350 23418 13356 23420
rect 13412 23418 13436 23420
rect 13492 23418 13516 23420
rect 13572 23418 13596 23420
rect 13652 23418 13658 23420
rect 13412 23366 13414 23418
rect 13594 23366 13596 23418
rect 13350 23364 13356 23366
rect 13412 23364 13436 23366
rect 13492 23364 13516 23366
rect 13572 23364 13596 23366
rect 13652 23364 13658 23366
rect 13350 23355 13658 23364
rect 13350 22332 13658 22341
rect 13350 22330 13356 22332
rect 13412 22330 13436 22332
rect 13492 22330 13516 22332
rect 13572 22330 13596 22332
rect 13652 22330 13658 22332
rect 13412 22278 13414 22330
rect 13594 22278 13596 22330
rect 13350 22276 13356 22278
rect 13412 22276 13436 22278
rect 13492 22276 13516 22278
rect 13572 22276 13596 22278
rect 13652 22276 13658 22278
rect 13350 22267 13658 22276
rect 13740 22166 13768 24210
rect 13832 24070 13860 24550
rect 14108 24206 14136 24550
rect 14200 24290 14228 26924
rect 14844 25242 14872 26924
rect 14752 25214 14872 25242
rect 14752 24818 14780 25214
rect 14850 25052 15158 25061
rect 14850 25050 14856 25052
rect 14912 25050 14936 25052
rect 14992 25050 15016 25052
rect 15072 25050 15096 25052
rect 15152 25050 15158 25052
rect 14912 24998 14914 25050
rect 15094 24998 15096 25050
rect 14850 24996 14856 24998
rect 14912 24996 14936 24998
rect 14992 24996 15016 24998
rect 15072 24996 15096 24998
rect 15152 24996 15158 24998
rect 14850 24987 15158 24996
rect 15488 24818 15516 26924
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14200 24262 14320 24290
rect 14292 24206 14320 24262
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 22642 13860 24006
rect 13924 23798 13952 24074
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 14094 23624 14150 23633
rect 14094 23559 14150 23568
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13556 21690 13584 21830
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13740 21486 13768 22102
rect 14004 21956 14056 21962
rect 14004 21898 14056 21904
rect 14016 21690 14044 21898
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13350 21244 13658 21253
rect 13350 21242 13356 21244
rect 13412 21242 13436 21244
rect 13492 21242 13516 21244
rect 13572 21242 13596 21244
rect 13652 21242 13658 21244
rect 13412 21190 13414 21242
rect 13594 21190 13596 21242
rect 13350 21188 13356 21190
rect 13412 21188 13436 21190
rect 13492 21188 13516 21190
rect 13572 21188 13596 21190
rect 13652 21188 13658 21190
rect 13350 21179 13658 21188
rect 13636 21072 13688 21078
rect 13634 21040 13636 21049
rect 13688 21040 13690 21049
rect 13634 20975 13690 20984
rect 13350 20156 13658 20165
rect 13350 20154 13356 20156
rect 13412 20154 13436 20156
rect 13492 20154 13516 20156
rect 13572 20154 13596 20156
rect 13652 20154 13658 20156
rect 13412 20102 13414 20154
rect 13594 20102 13596 20154
rect 13350 20100 13356 20102
rect 13412 20100 13436 20102
rect 13492 20100 13516 20102
rect 13572 20100 13596 20102
rect 13652 20100 13658 20102
rect 13350 20091 13658 20100
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13280 18766 13308 19450
rect 13740 19242 13768 21422
rect 14108 21146 14136 23559
rect 14200 22778 14228 24142
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14384 23050 14412 24006
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14200 21486 14228 22034
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13924 20058 13952 20878
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 14016 20466 14044 20742
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14108 19496 14136 21082
rect 14292 19904 14320 22374
rect 14384 22098 14412 22510
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14568 21978 14596 24006
rect 14660 23866 14688 24686
rect 14850 23964 15158 23973
rect 14850 23962 14856 23964
rect 14912 23962 14936 23964
rect 14992 23962 15016 23964
rect 15072 23962 15096 23964
rect 15152 23962 15158 23964
rect 14912 23910 14914 23962
rect 15094 23910 15096 23962
rect 14850 23908 14856 23910
rect 14912 23908 14936 23910
rect 14992 23908 15016 23910
rect 15072 23908 15096 23910
rect 15152 23908 15158 23910
rect 14850 23899 15158 23908
rect 14648 23860 14700 23866
rect 14700 23820 14872 23848
rect 14648 23802 14700 23808
rect 14844 23730 14872 23820
rect 14648 23724 14700 23730
rect 14832 23724 14884 23730
rect 14700 23684 14780 23712
rect 14648 23666 14700 23672
rect 14752 23322 14780 23684
rect 14832 23666 14884 23672
rect 15106 23624 15162 23633
rect 15106 23559 15108 23568
rect 15160 23559 15162 23568
rect 15108 23530 15160 23536
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14660 22778 14688 22986
rect 14850 22876 15158 22885
rect 14850 22874 14856 22876
rect 14912 22874 14936 22876
rect 14992 22874 15016 22876
rect 15072 22874 15096 22876
rect 15152 22874 15158 22876
rect 14912 22822 14914 22874
rect 15094 22822 15096 22874
rect 14850 22820 14856 22822
rect 14912 22820 14936 22822
rect 14992 22820 15016 22822
rect 15072 22820 15096 22822
rect 15152 22820 15158 22822
rect 14850 22811 15158 22820
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14660 22642 14688 22714
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14384 21950 14596 21978
rect 14384 21570 14412 21950
rect 14464 21888 14516 21894
rect 14660 21842 14688 22374
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14464 21830 14516 21836
rect 14476 21690 14504 21830
rect 14568 21814 14688 21842
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14384 21554 14504 21570
rect 14384 21548 14516 21554
rect 14384 21542 14464 21548
rect 14464 21490 14516 21496
rect 14476 20466 14504 21490
rect 14568 21350 14596 21814
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14556 21072 14608 21078
rect 14660 21060 14688 21626
rect 14608 21032 14688 21060
rect 14556 21014 14608 21020
rect 14752 20890 14780 21966
rect 14850 21788 15158 21797
rect 14850 21786 14856 21788
rect 14912 21786 14936 21788
rect 14992 21786 15016 21788
rect 15072 21786 15096 21788
rect 15152 21786 15158 21788
rect 14912 21734 14914 21786
rect 15094 21734 15096 21786
rect 14850 21732 14856 21734
rect 14912 21732 14936 21734
rect 14992 21732 15016 21734
rect 15072 21732 15096 21734
rect 15152 21732 15158 21734
rect 14850 21723 15158 21732
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15120 21049 15148 21082
rect 15106 21040 15162 21049
rect 15106 20975 15108 20984
rect 15160 20975 15162 20984
rect 15108 20946 15160 20952
rect 15016 20936 15068 20942
rect 14752 20884 15016 20890
rect 14752 20878 15068 20884
rect 14752 20862 15056 20878
rect 14752 20602 14780 20862
rect 14850 20700 15158 20709
rect 14850 20698 14856 20700
rect 14912 20698 14936 20700
rect 14992 20698 15016 20700
rect 15072 20698 15096 20700
rect 15152 20698 15158 20700
rect 14912 20646 14914 20698
rect 15094 20646 15096 20698
rect 14850 20644 14856 20646
rect 14912 20644 14936 20646
rect 14992 20644 15016 20646
rect 15072 20644 15096 20646
rect 15152 20644 15158 20646
rect 14850 20635 15158 20644
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 15212 20534 15240 23054
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14372 19916 14424 19922
rect 14292 19876 14372 19904
rect 14372 19858 14424 19864
rect 14108 19468 14320 19496
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13350 19068 13658 19077
rect 13350 19066 13356 19068
rect 13412 19066 13436 19068
rect 13492 19066 13516 19068
rect 13572 19066 13596 19068
rect 13652 19066 13658 19068
rect 13412 19014 13414 19066
rect 13594 19014 13596 19066
rect 13350 19012 13356 19014
rect 13412 19012 13436 19014
rect 13492 19012 13516 19014
rect 13572 19012 13596 19014
rect 13652 19012 13658 19014
rect 13350 19003 13658 19012
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13350 17980 13658 17989
rect 13350 17978 13356 17980
rect 13412 17978 13436 17980
rect 13492 17978 13516 17980
rect 13572 17978 13596 17980
rect 13652 17978 13658 17980
rect 13412 17926 13414 17978
rect 13594 17926 13596 17978
rect 13350 17924 13356 17926
rect 13412 17924 13436 17926
rect 13492 17924 13516 17926
rect 13572 17924 13596 17926
rect 13652 17924 13658 17926
rect 13350 17915 13658 17924
rect 13832 17542 13860 18770
rect 13924 18222 13952 19314
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 14200 17882 14228 19246
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14188 17672 14240 17678
rect 14292 17649 14320 19468
rect 14188 17614 14240 17620
rect 14278 17640 14334 17649
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13556 17270 13584 17478
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13350 16892 13658 16901
rect 13350 16890 13356 16892
rect 13412 16890 13436 16892
rect 13492 16890 13516 16892
rect 13572 16890 13596 16892
rect 13652 16890 13658 16892
rect 13412 16838 13414 16890
rect 13594 16838 13596 16890
rect 13350 16836 13356 16838
rect 13412 16836 13436 16838
rect 13492 16836 13516 16838
rect 13572 16836 13596 16838
rect 13652 16836 13658 16838
rect 13350 16827 13658 16836
rect 14108 16794 14136 17614
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 15162 12940 15302
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13004 15026 13032 15982
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13004 14634 13032 14962
rect 12912 14618 13032 14634
rect 12900 14612 13032 14618
rect 12952 14606 13032 14612
rect 12900 14554 12952 14560
rect 13096 14498 13124 15098
rect 13280 14958 13308 15914
rect 13350 15804 13658 15813
rect 13350 15802 13356 15804
rect 13412 15802 13436 15804
rect 13492 15802 13516 15804
rect 13572 15802 13596 15804
rect 13652 15802 13658 15804
rect 13412 15750 13414 15802
rect 13594 15750 13596 15802
rect 13350 15748 13356 15750
rect 13412 15748 13436 15750
rect 13492 15748 13516 15750
rect 13572 15748 13596 15750
rect 13652 15748 13658 15750
rect 13350 15739 13658 15748
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13924 14958 13952 15302
rect 14016 15162 14044 16050
rect 14200 15722 14228 17614
rect 14278 17575 14334 17584
rect 14384 16590 14412 19858
rect 14752 19854 14780 20402
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14850 19612 15158 19621
rect 14850 19610 14856 19612
rect 14912 19610 14936 19612
rect 14992 19610 15016 19612
rect 15072 19610 15096 19612
rect 15152 19610 15158 19612
rect 14912 19558 14914 19610
rect 15094 19558 15096 19610
rect 14850 19556 14856 19558
rect 14912 19556 14936 19558
rect 14992 19556 15016 19558
rect 15072 19556 15096 19558
rect 15152 19556 15158 19558
rect 14850 19547 15158 19556
rect 15304 19514 15332 24754
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23730 15608 24006
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15396 21146 15424 21966
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15488 21010 15516 23462
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15396 20602 15424 20742
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15396 19922 15424 20538
rect 15580 20398 15608 23122
rect 15672 22574 15700 23258
rect 15764 22982 15792 23598
rect 15856 23186 15884 23802
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15672 20602 15700 21830
rect 16040 21146 16068 24686
rect 16132 24614 16160 26924
rect 17850 25052 18158 25061
rect 17850 25050 17856 25052
rect 17912 25050 17936 25052
rect 17992 25050 18016 25052
rect 18072 25050 18096 25052
rect 18152 25050 18158 25052
rect 17912 24998 17914 25050
rect 18094 24998 18096 25050
rect 17850 24996 17856 24998
rect 17912 24996 17936 24998
rect 17992 24996 18016 24998
rect 18072 24996 18096 24998
rect 18152 24996 18158 24998
rect 17850 24987 18158 24996
rect 18708 24834 18736 26924
rect 18708 24818 18828 24834
rect 19352 24818 19380 26924
rect 19996 24818 20024 26924
rect 20850 25052 21158 25061
rect 20850 25050 20856 25052
rect 20912 25050 20936 25052
rect 20992 25050 21016 25052
rect 21072 25050 21096 25052
rect 21152 25050 21158 25052
rect 20912 24998 20914 25050
rect 21094 24998 21096 25050
rect 20850 24996 20856 24998
rect 20912 24996 20936 24998
rect 20992 24996 21016 24998
rect 21072 24996 21096 24998
rect 21152 24996 21158 24998
rect 20850 24987 21158 24996
rect 23850 25052 24158 25061
rect 23850 25050 23856 25052
rect 23912 25050 23936 25052
rect 23992 25050 24016 25052
rect 24072 25050 24096 25052
rect 24152 25050 24158 25052
rect 23912 24998 23914 25050
rect 24094 24998 24096 25050
rect 23850 24996 23856 24998
rect 23912 24996 23936 24998
rect 23992 24996 24016 24998
rect 24072 24996 24096 24998
rect 24152 24996 24158 24998
rect 23850 24987 24158 24996
rect 16212 24812 16264 24818
rect 18708 24812 18840 24818
rect 18708 24806 18788 24812
rect 16212 24754 16264 24760
rect 18788 24754 18840 24760
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16224 24410 16252 24754
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 16350 24508 16658 24517
rect 16350 24506 16356 24508
rect 16412 24506 16436 24508
rect 16492 24506 16516 24508
rect 16572 24506 16596 24508
rect 16652 24506 16658 24508
rect 16412 24454 16414 24506
rect 16594 24454 16596 24506
rect 16350 24452 16356 24454
rect 16412 24452 16436 24454
rect 16492 24452 16516 24454
rect 16572 24452 16596 24454
rect 16652 24452 16658 24454
rect 16350 24443 16658 24452
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 18236 24268 18288 24274
rect 18236 24210 18288 24216
rect 16224 23118 16252 24210
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16592 23866 16620 24074
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16350 23420 16658 23429
rect 16350 23418 16356 23420
rect 16412 23418 16436 23420
rect 16492 23418 16516 23420
rect 16572 23418 16596 23420
rect 16652 23418 16658 23420
rect 16412 23366 16414 23418
rect 16594 23366 16596 23418
rect 16350 23364 16356 23366
rect 16412 23364 16436 23366
rect 16492 23364 16516 23366
rect 16572 23364 16596 23366
rect 16652 23364 16658 23366
rect 16350 23355 16658 23364
rect 16776 23322 16804 23666
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22574 16436 22918
rect 16868 22778 16896 24074
rect 17850 23964 18158 23973
rect 17850 23962 17856 23964
rect 17912 23962 17936 23964
rect 17992 23962 18016 23964
rect 18072 23962 18096 23964
rect 18152 23962 18158 23964
rect 17912 23910 17914 23962
rect 18094 23910 18096 23962
rect 17850 23908 17856 23910
rect 17912 23908 17936 23910
rect 17992 23908 18016 23910
rect 18072 23908 18096 23910
rect 18152 23908 18158 23910
rect 17850 23899 18158 23908
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17144 22778 17172 22986
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17236 22642 17264 22986
rect 17328 22642 17356 23462
rect 17604 22778 17632 23598
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16350 22332 16658 22341
rect 16350 22330 16356 22332
rect 16412 22330 16436 22332
rect 16492 22330 16516 22332
rect 16572 22330 16596 22332
rect 16652 22330 16658 22332
rect 16412 22278 16414 22330
rect 16594 22278 16596 22330
rect 16350 22276 16356 22278
rect 16412 22276 16436 22278
rect 16492 22276 16516 22278
rect 16572 22276 16596 22278
rect 16652 22276 16658 22278
rect 16350 22267 16658 22276
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16316 21554 16344 21898
rect 16684 21690 16712 21966
rect 17696 21690 17724 23598
rect 18248 23118 18276 24210
rect 18340 23118 18368 24550
rect 18984 24138 19012 24550
rect 19076 24342 19104 24686
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18972 24132 19024 24138
rect 18972 24074 19024 24080
rect 18432 23662 18460 24074
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18786 23624 18842 23633
rect 18432 23186 18460 23598
rect 18616 23526 18644 23598
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18708 23322 18736 23598
rect 18786 23559 18842 23568
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18524 22930 18552 23122
rect 18432 22902 18552 22930
rect 17850 22876 18158 22885
rect 17850 22874 17856 22876
rect 17912 22874 17936 22876
rect 17992 22874 18016 22876
rect 18072 22874 18096 22876
rect 18152 22874 18158 22876
rect 17912 22822 17914 22874
rect 18094 22822 18096 22874
rect 17850 22820 17856 22822
rect 17912 22820 17936 22822
rect 17992 22820 18016 22822
rect 18072 22820 18096 22822
rect 18152 22820 18158 22822
rect 17850 22811 18158 22820
rect 18432 22166 18460 22902
rect 18708 22642 18736 23258
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 17850 21788 18158 21797
rect 17850 21786 17856 21788
rect 17912 21786 17936 21788
rect 17992 21786 18016 21788
rect 18072 21786 18096 21788
rect 18152 21786 18158 21788
rect 17912 21734 17914 21786
rect 18094 21734 18096 21786
rect 17850 21732 17856 21734
rect 17912 21732 17936 21734
rect 17992 21732 18016 21734
rect 18072 21732 18096 21734
rect 18152 21732 18158 21734
rect 17850 21723 18158 21732
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15856 20602 15884 20946
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14476 18426 14504 18702
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14660 18426 14688 18566
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14476 18290 14504 18362
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 17882 14596 18226
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14660 17762 14688 18362
rect 14476 17734 14688 17762
rect 14752 17762 14780 18566
rect 14850 18524 15158 18533
rect 14850 18522 14856 18524
rect 14912 18522 14936 18524
rect 14992 18522 15016 18524
rect 15072 18522 15096 18524
rect 15152 18522 15158 18524
rect 14912 18470 14914 18522
rect 15094 18470 15096 18522
rect 14850 18468 14856 18470
rect 14912 18468 14936 18470
rect 14992 18468 15016 18470
rect 15072 18468 15096 18470
rect 15152 18468 15158 18470
rect 14850 18459 15158 18468
rect 15304 18222 15332 18770
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15396 18426 15424 18702
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 14752 17734 14872 17762
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14476 16522 14504 17734
rect 14648 17672 14700 17678
rect 14554 17640 14610 17649
rect 14700 17632 14780 17660
rect 14648 17614 14700 17620
rect 14554 17575 14610 17584
rect 14568 17490 14596 17575
rect 14568 17462 14688 17490
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16658 14596 17002
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14660 16538 14688 17462
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14568 16510 14688 16538
rect 14108 15706 14228 15722
rect 14096 15700 14228 15706
rect 14148 15694 14228 15700
rect 14096 15642 14148 15648
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13004 14470 13124 14498
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 13004 13326 13032 14470
rect 13280 13530 13308 14894
rect 13350 14716 13658 14725
rect 13350 14714 13356 14716
rect 13412 14714 13436 14716
rect 13492 14714 13516 14716
rect 13572 14714 13596 14716
rect 13652 14714 13658 14716
rect 13412 14662 13414 14714
rect 13594 14662 13596 14714
rect 13350 14660 13356 14662
rect 13412 14660 13436 14662
rect 13492 14660 13516 14662
rect 13572 14660 13596 14662
rect 13652 14660 13658 14662
rect 13350 14651 13658 14660
rect 13740 14618 13768 14894
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13740 13977 13768 14010
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13350 13628 13658 13637
rect 13350 13626 13356 13628
rect 13412 13626 13436 13628
rect 13492 13626 13516 13628
rect 13572 13626 13596 13628
rect 13652 13626 13658 13628
rect 13412 13574 13414 13626
rect 13594 13574 13596 13626
rect 13350 13572 13356 13574
rect 13412 13572 13436 13574
rect 13492 13572 13516 13574
rect 13572 13572 13596 13574
rect 13652 13572 13658 13574
rect 13350 13563 13658 13572
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12636 12406 12756 12434
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 11850 11996 12158 12005
rect 11850 11994 11856 11996
rect 11912 11994 11936 11996
rect 11992 11994 12016 11996
rect 12072 11994 12096 11996
rect 12152 11994 12158 11996
rect 11912 11942 11914 11994
rect 12094 11942 12096 11994
rect 11850 11940 11856 11942
rect 11912 11940 11936 11942
rect 11992 11940 12016 11942
rect 12072 11940 12096 11942
rect 12152 11940 12158 11942
rect 11850 11931 12158 11940
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 12544 11218 12572 12038
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 11850 10908 12158 10917
rect 11850 10906 11856 10908
rect 11912 10906 11936 10908
rect 11992 10906 12016 10908
rect 12072 10906 12096 10908
rect 12152 10906 12158 10908
rect 11912 10854 11914 10906
rect 12094 10854 12096 10906
rect 11850 10852 11856 10854
rect 11912 10852 11936 10854
rect 11992 10852 12016 10854
rect 12072 10852 12096 10854
rect 12152 10852 12158 10854
rect 11850 10843 12158 10852
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11992 10266 12020 10678
rect 12636 10538 12664 12406
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 11850 9820 12158 9829
rect 11850 9818 11856 9820
rect 11912 9818 11936 9820
rect 11992 9818 12016 9820
rect 12072 9818 12096 9820
rect 12152 9818 12158 9820
rect 11912 9766 11914 9818
rect 12094 9766 12096 9818
rect 11850 9764 11856 9766
rect 11912 9764 11936 9766
rect 11992 9764 12016 9766
rect 12072 9764 12096 9766
rect 12152 9764 12158 9766
rect 11850 9755 12158 9764
rect 12452 9178 12480 9930
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9586 12572 9862
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12636 8974 12664 9318
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 7886 11560 8842
rect 12728 8786 12756 11698
rect 12636 8758 12756 8786
rect 11850 8732 12158 8741
rect 11850 8730 11856 8732
rect 11912 8730 11936 8732
rect 11992 8730 12016 8732
rect 12072 8730 12096 8732
rect 12152 8730 12158 8732
rect 11912 8678 11914 8730
rect 12094 8678 12096 8730
rect 11850 8676 11856 8678
rect 11912 8676 11936 8678
rect 11992 8676 12016 8678
rect 12072 8676 12096 8678
rect 12152 8676 12158 8678
rect 11850 8667 12158 8676
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11532 6746 11560 7822
rect 11716 7546 11744 8434
rect 12636 8022 12664 8758
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11850 7644 12158 7653
rect 11850 7642 11856 7644
rect 11912 7642 11936 7644
rect 11992 7642 12016 7644
rect 12072 7642 12096 7644
rect 12152 7642 12158 7644
rect 11912 7590 11914 7642
rect 12094 7590 12096 7642
rect 11850 7588 11856 7590
rect 11912 7588 11936 7590
rect 11992 7588 12016 7590
rect 12072 7588 12096 7590
rect 12152 7588 12158 7590
rect 11850 7579 12158 7588
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 12268 7410 12296 7686
rect 12636 7546 12664 7958
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12728 7478 12756 7754
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 6798 12480 7346
rect 12728 7002 12756 7414
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 11704 6792 11756 6798
rect 11532 6718 11652 6746
rect 11704 6734 11756 6740
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 8850 5468 9158 5477
rect 8850 5466 8856 5468
rect 8912 5466 8936 5468
rect 8992 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9158 5468
rect 8912 5414 8914 5466
rect 9094 5414 9096 5466
rect 8850 5412 8856 5414
rect 8912 5412 8936 5414
rect 8992 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9158 5414
rect 8850 5403 9158 5412
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8680 5234 8708 5306
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3126 8248 4014
rect 8312 3942 8340 4558
rect 8404 4146 8432 4558
rect 8588 4554 8616 5170
rect 8680 4690 8708 5170
rect 8864 4690 8892 5238
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8576 4548 8628 4554
rect 8864 4536 8892 4626
rect 8576 4490 8628 4496
rect 8680 4508 8892 4536
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8404 3738 8432 4082
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8496 3602 8524 4082
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8312 3398 8340 3538
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8312 2514 8340 3334
rect 8404 3194 8432 3470
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8588 2446 8616 4490
rect 8680 3670 8708 4508
rect 8956 4468 8984 5306
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 4758 9260 5102
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 8772 4440 8984 4468
rect 9220 4480 9272 4486
rect 8772 4010 8800 4440
rect 9220 4422 9272 4428
rect 8850 4380 9158 4389
rect 8850 4378 8856 4380
rect 8912 4378 8936 4380
rect 8992 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9158 4380
rect 8912 4326 8914 4378
rect 9094 4326 9096 4378
rect 8850 4324 8856 4326
rect 8912 4324 8936 4326
rect 8992 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9158 4326
rect 8850 4315 9158 4324
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 9232 3942 9260 4422
rect 9324 4010 9352 5646
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5098 9444 5510
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9588 4752 9640 4758
rect 9416 4700 9588 4706
rect 9416 4694 9640 4700
rect 9416 4678 9628 4694
rect 9416 4282 9444 4678
rect 9588 4616 9640 4622
rect 9508 4564 9588 4570
rect 9508 4558 9640 4564
rect 9508 4542 9628 4558
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9416 4146 9444 4218
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9508 4026 9536 4542
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9416 3998 9536 4026
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3738 9260 3878
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 9048 3466 9076 3674
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 9416 3398 9444 3998
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3670 9536 3878
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9600 3534 9628 4422
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9784 3670 9812 4014
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 8850 3292 9158 3301
rect 8850 3290 8856 3292
rect 8912 3290 8936 3292
rect 8992 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9158 3292
rect 8912 3238 8914 3290
rect 9094 3238 9096 3290
rect 8850 3236 8856 3238
rect 8912 3236 8936 3238
rect 8992 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9158 3238
rect 8850 3227 9158 3236
rect 9508 3194 9536 3402
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9508 2922 9536 3130
rect 9600 2990 9628 3470
rect 9784 3058 9812 3606
rect 9876 3466 9904 3946
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9968 2774 9996 5646
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 3058 10088 3334
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10152 2854 10180 6394
rect 11532 6390 11560 6598
rect 11624 6458 11652 6718
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 10350 6012 10658 6021
rect 10350 6010 10356 6012
rect 10412 6010 10436 6012
rect 10492 6010 10516 6012
rect 10572 6010 10596 6012
rect 10652 6010 10658 6012
rect 10412 5958 10414 6010
rect 10594 5958 10596 6010
rect 10350 5956 10356 5958
rect 10412 5956 10436 5958
rect 10492 5956 10516 5958
rect 10572 5956 10596 5958
rect 10652 5956 10658 5958
rect 10350 5947 10658 5956
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 10350 4924 10658 4933
rect 10350 4922 10356 4924
rect 10412 4922 10436 4924
rect 10492 4922 10516 4924
rect 10572 4922 10596 4924
rect 10652 4922 10658 4924
rect 10412 4870 10414 4922
rect 10594 4870 10596 4922
rect 10350 4868 10356 4870
rect 10412 4868 10436 4870
rect 10492 4868 10516 4870
rect 10572 4868 10596 4870
rect 10652 4868 10658 4870
rect 10350 4859 10658 4868
rect 11532 4826 11560 5578
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10244 3738 10272 4218
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10350 3836 10658 3845
rect 10350 3834 10356 3836
rect 10412 3834 10436 3836
rect 10492 3834 10516 3836
rect 10572 3834 10596 3836
rect 10652 3834 10658 3836
rect 10412 3782 10414 3834
rect 10594 3782 10596 3834
rect 10350 3780 10356 3782
rect 10412 3780 10436 3782
rect 10492 3780 10516 3782
rect 10572 3780 10596 3782
rect 10652 3780 10658 3782
rect 10350 3771 10658 3780
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10244 3466 10272 3674
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 10428 3194 10456 3538
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10704 3126 10732 4014
rect 10796 3738 10824 4422
rect 10888 4214 10916 4558
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10888 4010 10916 4150
rect 10980 4078 11008 4490
rect 11716 4146 11744 6734
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 11850 6556 12158 6565
rect 11850 6554 11856 6556
rect 11912 6554 11936 6556
rect 11992 6554 12016 6556
rect 12072 6554 12096 6556
rect 12152 6554 12158 6556
rect 11912 6502 11914 6554
rect 12094 6502 12096 6554
rect 11850 6500 11856 6502
rect 11912 6500 11936 6502
rect 11992 6500 12016 6502
rect 12072 6500 12096 6502
rect 12152 6500 12158 6502
rect 11850 6491 12158 6500
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 11850 5468 12158 5477
rect 11850 5466 11856 5468
rect 11912 5466 11936 5468
rect 11992 5466 12016 5468
rect 12072 5466 12096 5468
rect 12152 5466 12158 5468
rect 11912 5414 11914 5466
rect 12094 5414 12096 5466
rect 11850 5412 11856 5414
rect 11912 5412 11936 5414
rect 11992 5412 12016 5414
rect 12072 5412 12096 5414
rect 12152 5412 12158 5414
rect 11850 5403 12158 5412
rect 12268 4486 12296 6326
rect 12360 5914 12388 6598
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12452 5778 12480 6734
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4622 12388 4966
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 11850 4380 12158 4389
rect 11850 4378 11856 4380
rect 11912 4378 11936 4380
rect 11992 4378 12016 4380
rect 12072 4378 12096 4380
rect 12152 4378 12158 4380
rect 11912 4326 11914 4378
rect 12094 4326 12096 4378
rect 11850 4324 11856 4326
rect 11912 4324 11936 4326
rect 11992 4324 12016 4326
rect 12072 4324 12096 4326
rect 12152 4324 12158 4326
rect 11850 4315 12158 4324
rect 12268 4214 12296 4422
rect 12256 4208 12308 4214
rect 12176 4156 12256 4162
rect 12176 4150 12308 4156
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 12176 4134 12296 4150
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10796 3602 10824 3674
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10888 3482 10916 3946
rect 10796 3454 10916 3482
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10232 2984 10284 2990
rect 10284 2944 10456 2972
rect 10232 2926 10284 2932
rect 10428 2854 10456 2944
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 9692 2746 9996 2774
rect 10350 2748 10658 2757
rect 10350 2746 10356 2748
rect 10412 2746 10436 2748
rect 10492 2746 10516 2748
rect 10572 2746 10596 2748
rect 10652 2746 10658 2748
rect 9692 2514 9720 2746
rect 10412 2694 10414 2746
rect 10594 2694 10596 2746
rect 10350 2692 10356 2694
rect 10412 2692 10436 2694
rect 10492 2692 10516 2694
rect 10572 2692 10596 2694
rect 10652 2692 10658 2694
rect 10350 2683 10658 2692
rect 10796 2650 10824 3454
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 10888 2446 10916 3334
rect 10980 3058 11008 3334
rect 11348 3194 11376 4082
rect 12176 3466 12204 4134
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 11850 3292 12158 3301
rect 11850 3290 11856 3292
rect 11912 3290 11936 3292
rect 11992 3290 12016 3292
rect 12072 3290 12096 3292
rect 12152 3290 12158 3292
rect 11912 3238 11914 3290
rect 12094 3238 12096 3290
rect 11850 3236 11856 3238
rect 11912 3236 11936 3238
rect 11992 3236 12016 3238
rect 12072 3236 12096 3238
rect 12152 3236 12158 3238
rect 11850 3227 12158 3236
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 12452 2774 12480 5714
rect 12544 5642 12572 6666
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12452 2746 12572 2774
rect 12544 2582 12572 2746
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12820 2446 12848 12922
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12912 12238 12940 12718
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12912 11762 12940 12174
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12912 9586 12940 11698
rect 13004 11218 13032 12582
rect 13096 12102 13124 13466
rect 13176 13456 13228 13462
rect 13228 13404 13308 13410
rect 13176 13398 13308 13404
rect 13188 13382 13308 13398
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13096 11354 13124 11698
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 13004 10198 13032 10474
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13188 10062 13216 13194
rect 13280 12170 13308 13382
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13350 12540 13658 12549
rect 13350 12538 13356 12540
rect 13412 12538 13436 12540
rect 13492 12538 13516 12540
rect 13572 12538 13596 12540
rect 13652 12538 13658 12540
rect 13412 12486 13414 12538
rect 13594 12486 13596 12538
rect 13350 12484 13356 12486
rect 13412 12484 13436 12486
rect 13492 12484 13516 12486
rect 13572 12484 13596 12486
rect 13652 12484 13658 12486
rect 13350 12475 13658 12484
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13740 11558 13768 13330
rect 13832 11830 13860 14282
rect 13924 13938 13952 14894
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14108 12238 14136 15642
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14292 14482 14320 14758
rect 14476 14618 14504 14894
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14568 14550 14596 16510
rect 14752 15502 14780 17632
rect 14844 17610 14872 17734
rect 14936 17649 14964 18090
rect 15304 17882 15332 18158
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 14922 17640 14978 17649
rect 14832 17604 14884 17610
rect 14922 17575 14978 17584
rect 14832 17546 14884 17552
rect 14850 17436 15158 17445
rect 14850 17434 14856 17436
rect 14912 17434 14936 17436
rect 14992 17434 15016 17436
rect 15072 17434 15096 17436
rect 15152 17434 15158 17436
rect 14912 17382 14914 17434
rect 15094 17382 15096 17434
rect 14850 17380 14856 17382
rect 14912 17380 14936 17382
rect 14992 17380 15016 17382
rect 15072 17380 15096 17382
rect 15152 17380 15158 17382
rect 14850 17371 15158 17380
rect 15396 17338 15424 18158
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15396 17202 15424 17274
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 14850 16348 15158 16357
rect 14850 16346 14856 16348
rect 14912 16346 14936 16348
rect 14992 16346 15016 16348
rect 15072 16346 15096 16348
rect 15152 16346 15158 16348
rect 14912 16294 14914 16346
rect 15094 16294 15096 16346
rect 14850 16292 14856 16294
rect 14912 16292 14936 16294
rect 14992 16292 15016 16294
rect 15072 16292 15096 16294
rect 15152 16292 15158 16294
rect 14850 16283 15158 16292
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15120 15502 15148 15846
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 14752 15094 14780 15438
rect 14850 15260 15158 15269
rect 14850 15258 14856 15260
rect 14912 15258 14936 15260
rect 14992 15258 15016 15260
rect 15072 15258 15096 15260
rect 15152 15258 15158 15260
rect 14912 15206 14914 15258
rect 15094 15206 15096 15258
rect 14850 15204 14856 15206
rect 14912 15204 14936 15206
rect 14992 15204 15016 15206
rect 15072 15204 15096 15206
rect 15152 15204 15158 15206
rect 14850 15195 15158 15204
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14660 14346 14688 14894
rect 14648 14340 14700 14346
rect 15120 14328 15148 14962
rect 15120 14300 15240 14328
rect 14648 14282 14700 14288
rect 14850 14172 15158 14181
rect 14850 14170 14856 14172
rect 14912 14170 14936 14172
rect 14992 14170 15016 14172
rect 15072 14170 15096 14172
rect 15152 14170 15158 14172
rect 14912 14118 14914 14170
rect 15094 14118 15096 14170
rect 14850 14116 14856 14118
rect 14912 14116 14936 14118
rect 14992 14116 15016 14118
rect 15072 14116 15096 14118
rect 15152 14116 15158 14118
rect 14850 14107 15158 14116
rect 15212 14074 15240 14300
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15304 14006 15332 14214
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 13326 14412 13670
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 15304 13258 15332 13942
rect 15396 13938 15424 15846
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14752 12918 14780 13126
rect 14850 13084 15158 13093
rect 14850 13082 14856 13084
rect 14912 13082 14936 13084
rect 14992 13082 15016 13084
rect 15072 13082 15096 13084
rect 15152 13082 15158 13084
rect 14912 13030 14914 13082
rect 15094 13030 15096 13082
rect 14850 13028 14856 13030
rect 14912 13028 14936 13030
rect 14992 13028 15016 13030
rect 15072 13028 15096 13030
rect 15152 13028 15158 13030
rect 14850 13019 15158 13028
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12238 14504 12582
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14108 11898 14136 12174
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14850 11996 15158 12005
rect 14850 11994 14856 11996
rect 14912 11994 14936 11996
rect 14992 11994 15016 11996
rect 15072 11994 15096 11996
rect 15152 11994 15158 11996
rect 14912 11942 14914 11994
rect 15094 11942 15096 11994
rect 14850 11940 14856 11942
rect 14912 11940 14936 11942
rect 14992 11940 15016 11942
rect 15072 11940 15096 11942
rect 15152 11940 15158 11942
rect 14850 11931 15158 11940
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13350 11452 13658 11461
rect 13350 11450 13356 11452
rect 13412 11450 13436 11452
rect 13492 11450 13516 11452
rect 13572 11450 13596 11452
rect 13652 11450 13658 11452
rect 13412 11398 13414 11450
rect 13594 11398 13596 11450
rect 13350 11396 13356 11398
rect 13412 11396 13436 11398
rect 13492 11396 13516 11398
rect 13572 11396 13596 11398
rect 13652 11396 13658 11398
rect 13350 11387 13658 11396
rect 13740 11354 13768 11494
rect 13832 11354 13860 11766
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12912 9178 12940 9522
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13280 8090 13308 11086
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13350 10364 13658 10373
rect 13350 10362 13356 10364
rect 13412 10362 13436 10364
rect 13492 10362 13516 10364
rect 13572 10362 13596 10364
rect 13652 10362 13658 10364
rect 13412 10310 13414 10362
rect 13594 10310 13596 10362
rect 13350 10308 13356 10310
rect 13412 10308 13436 10310
rect 13492 10308 13516 10310
rect 13572 10308 13596 10310
rect 13652 10308 13658 10310
rect 13350 10299 13658 10308
rect 13740 10130 13952 10146
rect 13728 10124 13952 10130
rect 13780 10118 13952 10124
rect 13728 10066 13780 10072
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13350 9276 13658 9285
rect 13350 9274 13356 9276
rect 13412 9274 13436 9276
rect 13492 9274 13516 9276
rect 13572 9274 13596 9276
rect 13652 9274 13658 9276
rect 13412 9222 13414 9274
rect 13594 9222 13596 9274
rect 13350 9220 13356 9222
rect 13412 9220 13436 9222
rect 13492 9220 13516 9222
rect 13572 9220 13596 9222
rect 13652 9220 13658 9222
rect 13350 9211 13658 9220
rect 13832 8634 13860 9862
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13350 8188 13658 8197
rect 13350 8186 13356 8188
rect 13412 8186 13436 8188
rect 13492 8186 13516 8188
rect 13572 8186 13596 8188
rect 13652 8186 13658 8188
rect 13412 8134 13414 8186
rect 13594 8134 13596 8186
rect 13350 8132 13356 8134
rect 13412 8132 13436 8134
rect 13492 8132 13516 8134
rect 13572 8132 13596 8134
rect 13652 8132 13658 8134
rect 13350 8123 13658 8132
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7410 13216 7822
rect 13820 7744 13872 7750
rect 13924 7732 13952 10118
rect 14016 7886 14044 11018
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14108 10266 14136 10610
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14200 9994 14228 11698
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 11218 14320 11494
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14370 11112 14426 11121
rect 14280 11076 14332 11082
rect 14370 11047 14426 11056
rect 14280 11018 14332 11024
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14200 9518 14228 9930
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13872 7704 13952 7732
rect 13820 7686 13872 7692
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13188 6730 13216 7346
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13280 7002 13308 7142
rect 13350 7100 13658 7109
rect 13350 7098 13356 7100
rect 13412 7098 13436 7100
rect 13492 7098 13516 7100
rect 13572 7098 13596 7100
rect 13652 7098 13658 7100
rect 13412 7046 13414 7098
rect 13594 7046 13596 7098
rect 13350 7044 13356 7046
rect 13412 7044 13436 7046
rect 13492 7044 13516 7046
rect 13572 7044 13596 7046
rect 13652 7044 13658 7046
rect 13350 7035 13658 7044
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13280 6118 13308 6938
rect 13832 6934 13860 7686
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 14016 6730 14044 7822
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6322 13860 6598
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13280 5642 13308 6054
rect 13350 6012 13658 6021
rect 13350 6010 13356 6012
rect 13412 6010 13436 6012
rect 13492 6010 13516 6012
rect 13572 6010 13596 6012
rect 13652 6010 13658 6012
rect 13412 5958 13414 6010
rect 13594 5958 13596 6010
rect 13350 5956 13356 5958
rect 13412 5956 13436 5958
rect 13492 5956 13516 5958
rect 13572 5956 13596 5958
rect 13652 5956 13658 5958
rect 13350 5947 13658 5956
rect 14016 5710 14044 6054
rect 14108 5778 14136 6258
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13350 4924 13658 4933
rect 13350 4922 13356 4924
rect 13412 4922 13436 4924
rect 13492 4922 13516 4924
rect 13572 4922 13596 4924
rect 13652 4922 13658 4924
rect 13412 4870 13414 4922
rect 13594 4870 13596 4922
rect 13350 4868 13356 4870
rect 13412 4868 13436 4870
rect 13492 4868 13516 4870
rect 13572 4868 13596 4870
rect 13652 4868 13658 4870
rect 13350 4859 13658 4868
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 13004 2650 13032 4014
rect 13350 3836 13658 3845
rect 13350 3834 13356 3836
rect 13412 3834 13436 3836
rect 13492 3834 13516 3836
rect 13572 3834 13596 3836
rect 13652 3834 13658 3836
rect 13412 3782 13414 3834
rect 13594 3782 13596 3834
rect 13350 3780 13356 3782
rect 13412 3780 13436 3782
rect 13492 3780 13516 3782
rect 13572 3780 13596 3782
rect 13652 3780 13658 3782
rect 13350 3771 13658 3780
rect 13740 3738 13768 4082
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13832 3602 13860 4150
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 13188 3194 13216 3402
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13740 3058 13768 3334
rect 13832 3126 13860 3538
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14200 2774 14228 9454
rect 14292 7886 14320 11018
rect 14384 9586 14412 11047
rect 14850 10908 15158 10917
rect 14850 10906 14856 10908
rect 14912 10906 14936 10908
rect 14992 10906 15016 10908
rect 15072 10906 15096 10908
rect 15152 10906 15158 10908
rect 14912 10854 14914 10906
rect 15094 10854 15096 10906
rect 14850 10852 14856 10854
rect 14912 10852 14936 10854
rect 14992 10852 15016 10854
rect 15072 10852 15096 10854
rect 15152 10852 15158 10854
rect 14850 10843 15158 10852
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14384 8401 14412 9522
rect 14370 8392 14426 8401
rect 14370 8327 14426 8336
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7546 14320 7822
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14476 7426 14504 10406
rect 15028 10146 15056 10542
rect 15304 10198 15332 12038
rect 15488 11286 15516 17138
rect 15672 17066 15700 19178
rect 15856 18290 15884 20538
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19854 15976 20198
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16040 19156 16068 20334
rect 16132 20058 16160 21490
rect 16316 21434 16344 21490
rect 16224 21406 16344 21434
rect 16224 20534 16252 21406
rect 16350 21244 16658 21253
rect 16350 21242 16356 21244
rect 16412 21242 16436 21244
rect 16492 21242 16516 21244
rect 16572 21242 16596 21244
rect 16652 21242 16658 21244
rect 16412 21190 16414 21242
rect 16594 21190 16596 21242
rect 16350 21188 16356 21190
rect 16412 21188 16436 21190
rect 16492 21188 16516 21190
rect 16572 21188 16596 21190
rect 16652 21188 16658 21190
rect 16350 21179 16658 21188
rect 16868 21146 16896 21490
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 20534 16528 20878
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16224 19854 16252 20470
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16350 20156 16658 20165
rect 16350 20154 16356 20156
rect 16412 20154 16436 20156
rect 16492 20154 16516 20156
rect 16572 20154 16596 20156
rect 16652 20154 16658 20156
rect 16412 20102 16414 20154
rect 16594 20102 16596 20154
rect 16350 20100 16356 20102
rect 16412 20100 16436 20102
rect 16492 20100 16516 20102
rect 16572 20100 16596 20102
rect 16652 20100 16658 20102
rect 16350 20091 16658 20100
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16120 19168 16172 19174
rect 16040 19128 16120 19156
rect 16120 19110 16172 19116
rect 16132 18970 16160 19110
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18426 16068 18566
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16132 18222 16160 18906
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 16250 15976 16390
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16028 16176 16080 16182
rect 16224 16130 16252 19314
rect 16350 19068 16658 19077
rect 16350 19066 16356 19068
rect 16412 19066 16436 19068
rect 16492 19066 16516 19068
rect 16572 19066 16596 19068
rect 16652 19066 16658 19068
rect 16412 19014 16414 19066
rect 16594 19014 16596 19066
rect 16350 19012 16356 19014
rect 16412 19012 16436 19014
rect 16492 19012 16516 19014
rect 16572 19012 16596 19014
rect 16652 19012 16658 19014
rect 16350 19003 16658 19012
rect 16670 18320 16726 18329
rect 16776 18306 16804 20402
rect 16960 20330 16988 20810
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 17236 20058 17264 20334
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17696 19922 17724 21626
rect 18432 21010 18460 22102
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18524 20942 18552 21830
rect 18616 21690 18644 21830
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18696 21684 18748 21690
rect 18800 21672 18828 23559
rect 18892 22642 18920 24006
rect 19076 23662 19104 24278
rect 19168 24274 19196 24550
rect 19260 24410 19288 24686
rect 19350 24508 19658 24517
rect 19350 24506 19356 24508
rect 19412 24506 19436 24508
rect 19492 24506 19516 24508
rect 19572 24506 19596 24508
rect 19652 24506 19658 24508
rect 19412 24454 19414 24506
rect 19594 24454 19596 24506
rect 19350 24452 19356 24454
rect 19412 24452 19436 24454
rect 19492 24452 19516 24454
rect 19572 24452 19596 24454
rect 19652 24452 19658 24454
rect 19350 24443 19658 24452
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 19260 23662 19288 24346
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 19628 23798 19656 24074
rect 19616 23792 19668 23798
rect 19616 23734 19668 23740
rect 19064 23656 19116 23662
rect 19248 23656 19300 23662
rect 19064 23598 19116 23604
rect 19154 23624 19210 23633
rect 19248 23598 19300 23604
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19154 23559 19156 23568
rect 19208 23559 19210 23568
rect 19156 23530 19208 23536
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19350 23420 19658 23429
rect 19350 23418 19356 23420
rect 19412 23418 19436 23420
rect 19492 23418 19516 23420
rect 19572 23418 19596 23420
rect 19652 23418 19658 23420
rect 19412 23366 19414 23418
rect 19594 23366 19596 23418
rect 19350 23364 19356 23366
rect 19412 23364 19436 23366
rect 19492 23364 19516 23366
rect 19572 23364 19596 23366
rect 19652 23364 19658 23366
rect 19350 23355 19658 23364
rect 19904 23322 19932 23462
rect 19996 23322 20024 23598
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18984 21962 19012 23054
rect 19350 22332 19658 22341
rect 19350 22330 19356 22332
rect 19412 22330 19436 22332
rect 19492 22330 19516 22332
rect 19572 22330 19596 22332
rect 19652 22330 19658 22332
rect 19412 22278 19414 22330
rect 19594 22278 19596 22330
rect 19350 22276 19356 22278
rect 19412 22276 19436 22278
rect 19492 22276 19516 22278
rect 19572 22276 19596 22278
rect 19652 22276 19658 22278
rect 19350 22267 19658 22276
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18800 21644 18920 21672
rect 18696 21626 18748 21632
rect 18708 21570 18736 21626
rect 18616 21542 18736 21570
rect 18788 21548 18840 21554
rect 18616 21486 18644 21542
rect 18788 21490 18840 21496
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18800 21026 18828 21490
rect 18616 20998 18828 21026
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18616 20806 18644 20998
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 17850 20700 18158 20709
rect 17850 20698 17856 20700
rect 17912 20698 17936 20700
rect 17992 20698 18016 20700
rect 18072 20698 18096 20700
rect 18152 20698 18158 20700
rect 17912 20646 17914 20698
rect 18094 20646 18096 20698
rect 17850 20644 17856 20646
rect 17912 20644 17936 20646
rect 17992 20644 18016 20646
rect 18072 20644 18096 20646
rect 18152 20644 18158 20646
rect 17850 20635 18158 20644
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16726 18278 16804 18306
rect 16670 18255 16672 18264
rect 16724 18255 16726 18264
rect 16672 18226 16724 18232
rect 16350 17980 16658 17989
rect 16350 17978 16356 17980
rect 16412 17978 16436 17980
rect 16492 17978 16516 17980
rect 16572 17978 16596 17980
rect 16652 17978 16658 17980
rect 16412 17926 16414 17978
rect 16594 17926 16596 17978
rect 16350 17924 16356 17926
rect 16412 17924 16436 17926
rect 16492 17924 16516 17926
rect 16572 17924 16596 17926
rect 16652 17924 16658 17926
rect 16350 17915 16658 17924
rect 16868 17338 16896 18634
rect 16960 17610 16988 19450
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17420 18222 17448 18702
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16350 16892 16658 16901
rect 16350 16890 16356 16892
rect 16412 16890 16436 16892
rect 16492 16890 16516 16892
rect 16572 16890 16596 16892
rect 16652 16890 16658 16892
rect 16412 16838 16414 16890
rect 16594 16838 16596 16890
rect 16350 16836 16356 16838
rect 16412 16836 16436 16838
rect 16492 16836 16516 16838
rect 16572 16836 16596 16838
rect 16652 16836 16658 16838
rect 16350 16827 16658 16836
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16028 16118 16080 16124
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15580 14618 15608 16050
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 16040 14482 16068 16118
rect 16132 16114 16344 16130
rect 16132 16108 16356 16114
rect 16132 16102 16304 16108
rect 16132 15162 16160 16102
rect 16304 16050 16356 16056
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 14074 15884 14214
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 16132 13394 16160 14418
rect 16224 13462 16252 15982
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16350 15804 16658 15813
rect 16350 15802 16356 15804
rect 16412 15802 16436 15804
rect 16492 15802 16516 15804
rect 16572 15802 16596 15804
rect 16652 15802 16658 15804
rect 16412 15750 16414 15802
rect 16594 15750 16596 15802
rect 16350 15748 16356 15750
rect 16412 15748 16436 15750
rect 16492 15748 16516 15750
rect 16572 15748 16596 15750
rect 16652 15748 16658 15750
rect 16350 15739 16658 15748
rect 16776 15586 16804 15914
rect 16684 15570 16804 15586
rect 16672 15564 16804 15570
rect 16724 15558 16804 15564
rect 16672 15506 16724 15512
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15094 16528 15302
rect 16868 15162 16896 16526
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17215 15564 17267 15570
rect 17328 15552 17356 18090
rect 17420 17678 17448 18158
rect 17512 17814 17540 19858
rect 18616 19854 18644 20742
rect 18892 20058 18920 21644
rect 18984 21554 19012 21898
rect 19260 21554 19288 21966
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 18984 21162 19012 21490
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 18984 21134 19104 21162
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18984 20466 19012 21014
rect 19076 21010 19104 21134
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18984 19922 19012 20402
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 19168 19854 19196 21286
rect 19260 20398 19288 21490
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19350 21244 19658 21253
rect 19350 21242 19356 21244
rect 19412 21242 19436 21244
rect 19492 21242 19516 21244
rect 19572 21242 19596 21244
rect 19652 21242 19658 21244
rect 19412 21190 19414 21242
rect 19594 21190 19596 21242
rect 19350 21188 19356 21190
rect 19412 21188 19436 21190
rect 19492 21188 19516 21190
rect 19572 21188 19596 21190
rect 19652 21188 19658 21190
rect 19350 21179 19658 21188
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19352 20244 19380 20334
rect 19260 20216 19380 20244
rect 19260 20058 19288 20216
rect 19350 20156 19658 20165
rect 19350 20154 19356 20156
rect 19412 20154 19436 20156
rect 19492 20154 19516 20156
rect 19572 20154 19596 20156
rect 19652 20154 19658 20156
rect 19412 20102 19414 20154
rect 19594 20102 19596 20154
rect 19350 20100 19356 20102
rect 19412 20100 19436 20102
rect 19492 20100 19516 20102
rect 19572 20100 19596 20102
rect 19652 20100 19658 20102
rect 19350 20091 19658 20100
rect 19720 20058 19748 20810
rect 19812 20466 19840 21286
rect 19996 20602 20024 21490
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 17850 19612 18158 19621
rect 17850 19610 17856 19612
rect 17912 19610 17936 19612
rect 17992 19610 18016 19612
rect 18072 19610 18096 19612
rect 18152 19610 18158 19612
rect 17912 19558 17914 19610
rect 18094 19558 18096 19610
rect 17850 19556 17856 19558
rect 17912 19556 17936 19558
rect 17992 19556 18016 19558
rect 18072 19556 18096 19558
rect 18152 19556 18158 19558
rect 17850 19547 18158 19556
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17696 17882 17724 19314
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17420 17270 17448 17614
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17696 17202 17724 17614
rect 17788 17338 17816 19314
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 18604 18760 18656 18766
rect 18656 18720 18736 18748
rect 18604 18702 18656 18708
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 17850 18524 18158 18533
rect 17850 18522 17856 18524
rect 17912 18522 17936 18524
rect 17992 18522 18016 18524
rect 18072 18522 18096 18524
rect 18152 18522 18158 18524
rect 17912 18470 17914 18522
rect 18094 18470 18096 18522
rect 17850 18468 17856 18470
rect 17912 18468 17936 18470
rect 17992 18468 18016 18470
rect 18072 18468 18096 18470
rect 18152 18468 18158 18470
rect 17850 18459 18158 18468
rect 18248 17746 18276 18566
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18524 18222 18552 18362
rect 18708 18222 18736 18720
rect 18800 18698 18828 19246
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19350 19068 19658 19077
rect 19350 19066 19356 19068
rect 19412 19066 19436 19068
rect 19492 19066 19516 19068
rect 19572 19066 19596 19068
rect 19652 19066 19658 19068
rect 19412 19014 19414 19066
rect 19594 19014 19596 19066
rect 19350 19012 19356 19014
rect 19412 19012 19436 19014
rect 19492 19012 19516 19014
rect 19572 19012 19596 19014
rect 19652 19012 19658 19014
rect 19350 19003 19658 19012
rect 19720 18834 19748 19110
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 18788 18692 18840 18698
rect 18788 18634 18840 18640
rect 18800 18290 18828 18634
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 17850 17436 18158 17445
rect 17850 17434 17856 17436
rect 17912 17434 17936 17436
rect 17992 17434 18016 17436
rect 18072 17434 18096 17436
rect 18152 17434 18158 17436
rect 17912 17382 17914 17434
rect 18094 17382 18096 17434
rect 17850 17380 17856 17382
rect 17912 17380 17936 17382
rect 17992 17380 18016 17382
rect 18072 17380 18096 17382
rect 18152 17380 18158 17382
rect 17850 17371 18158 17380
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 15978 17724 16526
rect 18524 16522 18552 17614
rect 18708 17610 18736 18158
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17270 18644 17478
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18800 16794 18828 17614
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 19076 16658 19104 17002
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 17850 16348 18158 16357
rect 17850 16346 17856 16348
rect 17912 16346 17936 16348
rect 17992 16346 18016 16348
rect 18072 16346 18096 16348
rect 18152 16346 18158 16348
rect 17912 16294 17914 16346
rect 18094 16294 18096 16346
rect 17850 16292 17856 16294
rect 17912 16292 17936 16294
rect 17992 16292 18016 16294
rect 18072 16292 18096 16294
rect 18152 16292 18158 16294
rect 17850 16283 18158 16292
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17512 15570 17540 15642
rect 17267 15524 17356 15552
rect 17215 15506 17267 15512
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16350 14716 16658 14725
rect 16350 14714 16356 14716
rect 16412 14714 16436 14716
rect 16492 14714 16516 14716
rect 16572 14714 16596 14716
rect 16652 14714 16658 14716
rect 16412 14662 16414 14714
rect 16594 14662 16596 14714
rect 16350 14660 16356 14662
rect 16412 14660 16436 14662
rect 16492 14660 16516 14662
rect 16572 14660 16596 14662
rect 16652 14660 16658 14662
rect 16350 14651 16658 14660
rect 16960 14550 16988 14894
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 17052 14482 17080 15506
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 17236 14414 17264 14758
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 16350 13628 16658 13637
rect 16350 13626 16356 13628
rect 16412 13626 16436 13628
rect 16492 13626 16516 13628
rect 16572 13626 16596 13628
rect 16652 13626 16658 13628
rect 16412 13574 16414 13626
rect 16594 13574 16596 13626
rect 16350 13572 16356 13574
rect 16412 13572 16436 13574
rect 16492 13572 16516 13574
rect 16572 13572 16596 13574
rect 16652 13572 16658 13574
rect 16350 13563 16658 13572
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12170 15884 13126
rect 15948 12986 15976 13262
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16040 12442 16068 12854
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15672 11082 15700 11494
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 14568 10130 15056 10146
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 14568 10124 15068 10130
rect 14568 10118 15016 10124
rect 14568 9722 14596 10118
rect 15016 10066 15068 10072
rect 14832 10056 14884 10062
rect 14660 10016 14832 10044
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14568 8430 14596 9386
rect 14660 8838 14688 10016
rect 14832 9998 14884 10004
rect 14850 9820 15158 9829
rect 14850 9818 14856 9820
rect 14912 9818 14936 9820
rect 14992 9818 15016 9820
rect 15072 9818 15096 9820
rect 15152 9818 15158 9820
rect 14912 9766 14914 9818
rect 15094 9766 15096 9818
rect 14850 9764 14856 9766
rect 14912 9764 14936 9766
rect 14992 9764 15016 9766
rect 15072 9764 15096 9766
rect 15152 9764 15158 9766
rect 14850 9755 15158 9764
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15212 9178 15240 9454
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15212 9042 15240 9114
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8498 14688 8774
rect 14752 8634 14780 8842
rect 14850 8732 15158 8741
rect 14850 8730 14856 8732
rect 14912 8730 14936 8732
rect 14992 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15158 8732
rect 14912 8678 14914 8730
rect 15094 8678 15096 8730
rect 14850 8676 14856 8678
rect 14912 8676 14936 8678
rect 14992 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15158 8678
rect 14850 8667 15158 8676
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 15212 8566 15240 8978
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15304 8498 15332 9318
rect 15672 8974 15700 11018
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 9722 15792 10406
rect 15856 10130 15884 10542
rect 15948 10130 15976 11562
rect 16132 11558 16160 13330
rect 16224 12306 16252 13398
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16350 12540 16658 12549
rect 16350 12538 16356 12540
rect 16412 12538 16436 12540
rect 16492 12538 16516 12540
rect 16572 12538 16596 12540
rect 16652 12538 16658 12540
rect 16412 12486 16414 12538
rect 16594 12486 16596 12538
rect 16350 12484 16356 12486
rect 16412 12484 16436 12486
rect 16492 12484 16516 12486
rect 16572 12484 16596 12486
rect 16652 12484 16658 12486
rect 16350 12475 16658 12484
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11898 16528 12038
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16592 11762 16620 12378
rect 17144 12238 17172 13126
rect 17328 12782 17356 15524
rect 17500 15564 17552 15570
rect 17408 15512 17460 15518
rect 17500 15506 17552 15512
rect 17408 15454 17460 15460
rect 17420 15162 17448 15454
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16868 11762 16896 12174
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11354 16160 11494
rect 16350 11452 16658 11461
rect 16350 11450 16356 11452
rect 16412 11450 16436 11452
rect 16492 11450 16516 11452
rect 16572 11450 16596 11452
rect 16652 11450 16658 11452
rect 16412 11398 16414 11450
rect 16594 11398 16596 11450
rect 16350 11396 16356 11398
rect 16412 11396 16436 11398
rect 16492 11396 16516 11398
rect 16572 11396 16596 11398
rect 16652 11396 16658 11398
rect 16350 11387 16658 11396
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16408 10742 16436 11018
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 10248 16252 10406
rect 16350 10364 16658 10373
rect 16350 10362 16356 10364
rect 16412 10362 16436 10364
rect 16492 10362 16516 10364
rect 16572 10362 16596 10364
rect 16652 10362 16658 10364
rect 16412 10310 16414 10362
rect 16594 10310 16596 10362
rect 16350 10308 16356 10310
rect 16412 10308 16436 10310
rect 16492 10308 16516 10310
rect 16572 10308 16596 10310
rect 16652 10308 16658 10310
rect 16350 10299 16658 10308
rect 16224 10220 16344 10248
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15856 9178 15884 10066
rect 16120 10056 16172 10062
rect 16040 10016 16120 10044
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 16040 9042 16068 10016
rect 16120 9998 16172 10004
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16224 9178 16252 9862
rect 16316 9450 16344 10220
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16684 9722 16712 9930
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16350 9276 16658 9285
rect 16350 9274 16356 9276
rect 16412 9274 16436 9276
rect 16492 9274 16516 9276
rect 16572 9274 16596 9276
rect 16652 9274 16658 9276
rect 16412 9222 16414 9274
rect 16594 9222 16596 9274
rect 16350 9220 16356 9222
rect 16412 9220 16436 9222
rect 16492 9220 16516 9222
rect 16572 9220 16596 9222
rect 16652 9220 16658 9222
rect 16350 9211 16658 9220
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16316 8634 16344 8842
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7750 14596 8366
rect 16592 8362 16620 8774
rect 16776 8634 16804 9522
rect 16868 8974 16896 11698
rect 17328 11286 17356 12718
rect 17420 11830 17448 13126
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17512 11354 17540 13262
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12850 17632 13126
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17696 12238 17724 15914
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17788 13802 17816 15574
rect 18616 15570 18644 15982
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17850 15260 18158 15269
rect 17850 15258 17856 15260
rect 17912 15258 17936 15260
rect 17992 15258 18016 15260
rect 18072 15258 18096 15260
rect 18152 15258 18158 15260
rect 17912 15206 17914 15258
rect 18094 15206 18096 15258
rect 17850 15204 17856 15206
rect 17912 15204 17936 15206
rect 17992 15204 18016 15206
rect 18072 15204 18096 15206
rect 18152 15204 18158 15206
rect 17850 15195 18158 15204
rect 18248 14618 18276 15438
rect 18616 15162 18644 15506
rect 18800 15366 18828 16118
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18800 15162 18828 15302
rect 18984 15162 19012 15846
rect 19168 15620 19196 18090
rect 19352 18068 19380 18702
rect 19708 18352 19760 18358
rect 19812 18340 19840 19246
rect 19892 19236 19944 19242
rect 19892 19178 19944 19184
rect 19904 18766 19932 19178
rect 20180 18834 20208 24074
rect 20272 22778 20300 24074
rect 20456 23866 20484 24754
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20364 21146 20392 21966
rect 20456 21690 20484 23598
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20364 20602 20392 21082
rect 20732 20942 20760 24550
rect 22350 24508 22658 24517
rect 22350 24506 22356 24508
rect 22412 24506 22436 24508
rect 22492 24506 22516 24508
rect 22572 24506 22596 24508
rect 22652 24506 22658 24508
rect 22412 24454 22414 24506
rect 22594 24454 22596 24506
rect 22350 24452 22356 24454
rect 22412 24452 22436 24454
rect 22492 24452 22516 24454
rect 22572 24452 22596 24454
rect 22652 24452 22658 24454
rect 22350 24443 22658 24452
rect 20850 23964 21158 23973
rect 20850 23962 20856 23964
rect 20912 23962 20936 23964
rect 20992 23962 21016 23964
rect 21072 23962 21096 23964
rect 21152 23962 21158 23964
rect 20912 23910 20914 23962
rect 21094 23910 21096 23962
rect 20850 23908 20856 23910
rect 20912 23908 20936 23910
rect 20992 23908 21016 23910
rect 21072 23908 21096 23910
rect 21152 23908 21158 23910
rect 20850 23899 21158 23908
rect 23850 23964 24158 23973
rect 23850 23962 23856 23964
rect 23912 23962 23936 23964
rect 23992 23962 24016 23964
rect 24072 23962 24096 23964
rect 24152 23962 24158 23964
rect 23912 23910 23914 23962
rect 24094 23910 24096 23962
rect 23850 23908 23856 23910
rect 23912 23908 23936 23910
rect 23992 23908 24016 23910
rect 24072 23908 24096 23910
rect 24152 23908 24158 23910
rect 23850 23899 24158 23908
rect 22350 23420 22658 23429
rect 22350 23418 22356 23420
rect 22412 23418 22436 23420
rect 22492 23418 22516 23420
rect 22572 23418 22596 23420
rect 22652 23418 22658 23420
rect 22412 23366 22414 23418
rect 22594 23366 22596 23418
rect 22350 23364 22356 23366
rect 22412 23364 22436 23366
rect 22492 23364 22516 23366
rect 22572 23364 22596 23366
rect 22652 23364 22658 23366
rect 22350 23355 22658 23364
rect 20850 22876 21158 22885
rect 20850 22874 20856 22876
rect 20912 22874 20936 22876
rect 20992 22874 21016 22876
rect 21072 22874 21096 22876
rect 21152 22874 21158 22876
rect 20912 22822 20914 22874
rect 21094 22822 21096 22874
rect 20850 22820 20856 22822
rect 20912 22820 20936 22822
rect 20992 22820 21016 22822
rect 21072 22820 21096 22822
rect 21152 22820 21158 22822
rect 20850 22811 21158 22820
rect 23850 22876 24158 22885
rect 23850 22874 23856 22876
rect 23912 22874 23936 22876
rect 23992 22874 24016 22876
rect 24072 22874 24096 22876
rect 24152 22874 24158 22876
rect 23912 22822 23914 22874
rect 24094 22822 24096 22874
rect 23850 22820 23856 22822
rect 23912 22820 23936 22822
rect 23992 22820 24016 22822
rect 24072 22820 24096 22822
rect 24152 22820 24158 22822
rect 23850 22811 24158 22820
rect 22350 22332 22658 22341
rect 22350 22330 22356 22332
rect 22412 22330 22436 22332
rect 22492 22330 22516 22332
rect 22572 22330 22596 22332
rect 22652 22330 22658 22332
rect 22412 22278 22414 22330
rect 22594 22278 22596 22330
rect 22350 22276 22356 22278
rect 22412 22276 22436 22278
rect 22492 22276 22516 22278
rect 22572 22276 22596 22278
rect 22652 22276 22658 22278
rect 22350 22267 22658 22276
rect 20850 21788 21158 21797
rect 20850 21786 20856 21788
rect 20912 21786 20936 21788
rect 20992 21786 21016 21788
rect 21072 21786 21096 21788
rect 21152 21786 21158 21788
rect 20912 21734 20914 21786
rect 21094 21734 21096 21786
rect 20850 21732 20856 21734
rect 20912 21732 20936 21734
rect 20992 21732 21016 21734
rect 21072 21732 21096 21734
rect 21152 21732 21158 21734
rect 20850 21723 21158 21732
rect 23850 21788 24158 21797
rect 23850 21786 23856 21788
rect 23912 21786 23936 21788
rect 23992 21786 24016 21788
rect 24072 21786 24096 21788
rect 24152 21786 24158 21788
rect 23912 21734 23914 21786
rect 24094 21734 24096 21786
rect 23850 21732 23856 21734
rect 23912 21732 23936 21734
rect 23992 21732 24016 21734
rect 24072 21732 24096 21734
rect 24152 21732 24158 21734
rect 23850 21723 24158 21732
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 21010 21220 21286
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20732 20534 20760 20742
rect 20850 20700 21158 20709
rect 20850 20698 20856 20700
rect 20912 20698 20936 20700
rect 20992 20698 21016 20700
rect 21072 20698 21096 20700
rect 21152 20698 21158 20700
rect 20912 20646 20914 20698
rect 21094 20646 21096 20698
rect 20850 20644 20856 20646
rect 20912 20644 20936 20646
rect 20992 20644 21016 20646
rect 21072 20644 21096 20646
rect 21152 20644 21158 20646
rect 20850 20635 21158 20644
rect 21284 20602 21312 21490
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 22350 21244 22658 21253
rect 22350 21242 22356 21244
rect 22412 21242 22436 21244
rect 22492 21242 22516 21244
rect 22572 21242 22596 21244
rect 22652 21242 22658 21244
rect 22412 21190 22414 21242
rect 22594 21190 22596 21242
rect 22350 21188 22356 21190
rect 22412 21188 22436 21190
rect 22492 21188 22516 21190
rect 22572 21188 22596 21190
rect 22652 21188 22658 21190
rect 22350 21179 22658 21188
rect 23584 21185 23612 21286
rect 23570 21176 23626 21185
rect 23570 21111 23626 21120
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20850 19612 21158 19621
rect 20850 19610 20856 19612
rect 20912 19610 20936 19612
rect 20992 19610 21016 19612
rect 21072 19610 21096 19612
rect 21152 19610 21158 19612
rect 20912 19558 20914 19610
rect 21094 19558 21096 19610
rect 20850 19556 20856 19558
rect 20912 19556 20936 19558
rect 20992 19556 21016 19558
rect 21072 19556 21096 19558
rect 21152 19556 21158 19558
rect 20850 19547 21158 19556
rect 20720 19372 20772 19378
rect 20548 19320 20720 19334
rect 20548 19314 20772 19320
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20548 19306 20760 19314
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19996 18426 20024 18634
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19760 18312 19840 18340
rect 19708 18294 19760 18300
rect 19260 18040 19380 18068
rect 19260 17746 19288 18040
rect 19350 17980 19658 17989
rect 19350 17978 19356 17980
rect 19412 17978 19436 17980
rect 19492 17978 19516 17980
rect 19572 17978 19596 17980
rect 19652 17978 19658 17980
rect 19412 17926 19414 17978
rect 19594 17926 19596 17978
rect 19350 17924 19356 17926
rect 19412 17924 19436 17926
rect 19492 17924 19516 17926
rect 19572 17924 19596 17926
rect 19652 17924 19658 17926
rect 19350 17915 19658 17924
rect 19720 17882 19748 18294
rect 20180 18290 20208 18770
rect 20456 18766 20484 19110
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19904 17338 19932 18158
rect 20180 17610 20208 18226
rect 20272 17610 20300 18566
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20364 17338 20392 18226
rect 20548 17626 20576 19306
rect 20850 18524 21158 18533
rect 20850 18522 20856 18524
rect 20912 18522 20936 18524
rect 20992 18522 21016 18524
rect 21072 18522 21096 18524
rect 21152 18522 21158 18524
rect 20912 18470 20914 18522
rect 21094 18470 21096 18522
rect 20850 18468 20856 18470
rect 20912 18468 20936 18470
rect 20992 18468 21016 18470
rect 21072 18468 21096 18470
rect 21152 18468 21158 18470
rect 20850 18459 21158 18468
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20456 17598 20576 17626
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 19350 16892 19658 16901
rect 19350 16890 19356 16892
rect 19412 16890 19436 16892
rect 19492 16890 19516 16892
rect 19572 16890 19596 16892
rect 19652 16890 19658 16892
rect 19412 16838 19414 16890
rect 19594 16838 19596 16890
rect 19350 16836 19356 16838
rect 19412 16836 19436 16838
rect 19492 16836 19516 16838
rect 19572 16836 19596 16838
rect 19652 16836 19658 16838
rect 19350 16827 19658 16836
rect 20456 16794 20484 17598
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20548 17202 20576 17478
rect 20640 17270 20668 17614
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20640 16590 20668 17206
rect 20732 17202 20760 17847
rect 20850 17436 21158 17445
rect 20850 17434 20856 17436
rect 20912 17434 20936 17436
rect 20992 17434 21016 17436
rect 21072 17434 21096 17436
rect 21152 17434 21158 17436
rect 20912 17382 20914 17434
rect 21094 17382 21096 17434
rect 20850 17380 20856 17382
rect 20912 17380 20936 17382
rect 20992 17380 21016 17382
rect 21072 17380 21096 17382
rect 21152 17380 21158 17382
rect 20850 17371 21158 17380
rect 21284 17320 21312 19314
rect 21376 18970 21404 20946
rect 23850 20700 24158 20709
rect 23850 20698 23856 20700
rect 23912 20698 23936 20700
rect 23992 20698 24016 20700
rect 24072 20698 24096 20700
rect 24152 20698 24158 20700
rect 23912 20646 23914 20698
rect 24094 20646 24096 20698
rect 23850 20644 23856 20646
rect 23912 20644 23936 20646
rect 23992 20644 24016 20646
rect 24072 20644 24096 20646
rect 24152 20644 24158 20646
rect 23850 20635 24158 20644
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21100 17292 21312 17320
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 15910 20668 16186
rect 20732 16182 20760 17138
rect 21100 16590 21128 17292
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20850 16348 21158 16357
rect 20850 16346 20856 16348
rect 20912 16346 20936 16348
rect 20992 16346 21016 16348
rect 21072 16346 21096 16348
rect 21152 16346 21158 16348
rect 20912 16294 20914 16346
rect 21094 16294 21096 16346
rect 20850 16292 20856 16294
rect 20912 16292 20936 16294
rect 20992 16292 21016 16294
rect 21072 16292 21096 16294
rect 21152 16292 21158 16294
rect 20850 16283 21158 16292
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 19350 15804 19658 15813
rect 19350 15802 19356 15804
rect 19412 15802 19436 15804
rect 19492 15802 19516 15804
rect 19572 15802 19596 15804
rect 19652 15802 19658 15804
rect 19412 15750 19414 15802
rect 19594 15750 19596 15802
rect 19350 15748 19356 15750
rect 19412 15748 19436 15750
rect 19492 15748 19516 15750
rect 19572 15748 19596 15750
rect 19652 15748 19658 15750
rect 19350 15739 19658 15748
rect 19248 15632 19300 15638
rect 19168 15600 19248 15620
rect 19300 15600 19302 15609
rect 19168 15592 19246 15600
rect 19246 15535 19302 15544
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18984 14958 19012 15098
rect 19352 14958 19380 15438
rect 19812 15434 19840 15846
rect 20640 15586 20668 15846
rect 20732 15706 20760 15982
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20640 15558 20760 15586
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18972 14952 19024 14958
rect 19340 14952 19392 14958
rect 18972 14894 19024 14900
rect 19260 14900 19340 14906
rect 19260 14894 19392 14900
rect 18892 14618 18920 14894
rect 19260 14878 19380 14894
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 17850 14172 18158 14181
rect 17850 14170 17856 14172
rect 17912 14170 17936 14172
rect 17992 14170 18016 14172
rect 18072 14170 18096 14172
rect 18152 14170 18158 14172
rect 17912 14118 17914 14170
rect 18094 14118 18096 14170
rect 17850 14116 17856 14118
rect 17912 14116 17936 14118
rect 17992 14116 18016 14118
rect 18072 14116 18096 14118
rect 18152 14116 18158 14118
rect 17850 14107 18158 14116
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17788 12866 17816 13738
rect 19260 13716 19288 14878
rect 19350 14716 19658 14725
rect 19350 14714 19356 14716
rect 19412 14714 19436 14716
rect 19492 14714 19516 14716
rect 19572 14714 19596 14716
rect 19652 14714 19658 14716
rect 19412 14662 19414 14714
rect 19594 14662 19596 14714
rect 19350 14660 19356 14662
rect 19412 14660 19436 14662
rect 19492 14660 19516 14662
rect 19572 14660 19596 14662
rect 19652 14660 19658 14662
rect 19350 14651 19658 14660
rect 19996 14618 20024 14962
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19168 13688 19288 13716
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 17850 13084 18158 13093
rect 17850 13082 17856 13084
rect 17912 13082 17936 13084
rect 17992 13082 18016 13084
rect 18072 13082 18096 13084
rect 18152 13082 18158 13084
rect 17912 13030 17914 13082
rect 18094 13030 18096 13082
rect 17850 13028 17856 13030
rect 17912 13028 17936 13030
rect 17992 13028 18016 13030
rect 18072 13028 18096 13030
rect 18152 13028 18158 13030
rect 17850 13019 18158 13028
rect 17788 12838 17908 12866
rect 17880 12782 17908 12838
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 17788 12442 17816 12718
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11898 17724 12174
rect 18248 12102 18276 12650
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17850 11996 18158 12005
rect 17850 11994 17856 11996
rect 17912 11994 17936 11996
rect 17992 11994 18016 11996
rect 18072 11994 18096 11996
rect 18152 11994 18158 11996
rect 17912 11942 17914 11994
rect 18094 11942 18096 11994
rect 17850 11940 17856 11942
rect 17912 11940 17936 11942
rect 17992 11940 18016 11942
rect 18072 11940 18096 11942
rect 18152 11940 18158 11942
rect 17850 11931 18158 11940
rect 18340 11898 18368 12718
rect 18432 12442 18460 13330
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18800 12986 18828 13194
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 19168 12918 19196 13688
rect 19350 13628 19658 13637
rect 19350 13626 19356 13628
rect 19412 13626 19436 13628
rect 19492 13626 19516 13628
rect 19572 13626 19596 13628
rect 19652 13626 19658 13628
rect 19412 13574 19414 13626
rect 19594 13574 19596 13626
rect 19350 13572 19356 13574
rect 19412 13572 19436 13574
rect 19492 13572 19516 13574
rect 19572 13572 19596 13574
rect 19652 13572 19658 13574
rect 19350 13563 19658 13572
rect 20456 13410 20484 15098
rect 20732 15026 20760 15558
rect 20824 15502 20852 15846
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 21100 15434 21128 16050
rect 21192 15978 21220 16594
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 21284 15706 21312 17138
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20850 15260 21158 15269
rect 20850 15258 20856 15260
rect 20912 15258 20936 15260
rect 20992 15258 21016 15260
rect 21072 15258 21096 15260
rect 21152 15258 21158 15260
rect 20912 15206 20914 15258
rect 21094 15206 21096 15258
rect 20850 15204 20856 15206
rect 20912 15204 20936 15206
rect 20992 15204 21016 15206
rect 21072 15204 21096 15206
rect 21152 15204 21158 15206
rect 20850 15195 21158 15204
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 13954 20760 14962
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20824 14414 20852 14758
rect 21008 14618 21036 14894
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 21376 14226 21404 15914
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21468 14346 21496 15302
rect 21546 15056 21602 15065
rect 21546 14991 21602 15000
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21376 14198 21496 14226
rect 20850 14172 21158 14181
rect 20850 14170 20856 14172
rect 20912 14170 20936 14172
rect 20992 14170 21016 14172
rect 21072 14170 21096 14172
rect 21152 14170 21158 14172
rect 20912 14118 20914 14170
rect 21094 14118 21096 14170
rect 20850 14116 20856 14118
rect 20912 14116 20936 14118
rect 20992 14116 21016 14118
rect 21072 14116 21096 14118
rect 21152 14116 21158 14118
rect 20850 14107 21158 14116
rect 20812 14000 20864 14006
rect 20732 13948 20812 13954
rect 20732 13942 20864 13948
rect 20732 13926 20852 13942
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20456 13394 20668 13410
rect 20456 13388 20680 13394
rect 20456 13382 20628 13388
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19168 12782 19196 12854
rect 19444 12850 19472 13126
rect 19904 12986 19932 13126
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 20272 12782 20300 13126
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 19168 12306 19196 12718
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19350 12540 19658 12549
rect 19350 12538 19356 12540
rect 19412 12538 19436 12540
rect 19492 12538 19516 12540
rect 19572 12538 19596 12540
rect 19652 12538 19658 12540
rect 19412 12486 19414 12538
rect 19594 12486 19596 12538
rect 19350 12484 19356 12486
rect 19412 12484 19436 12486
rect 19492 12484 19516 12486
rect 19572 12484 19596 12486
rect 19652 12484 19658 12486
rect 19350 12475 19658 12484
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19812 12238 19840 12582
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 18340 11218 18368 11834
rect 18616 11762 18644 12038
rect 18708 11830 18736 12038
rect 19260 11898 19288 12038
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18708 11354 18736 11766
rect 19350 11452 19658 11461
rect 19350 11450 19356 11452
rect 19412 11450 19436 11452
rect 19492 11450 19516 11452
rect 19572 11450 19596 11452
rect 19652 11450 19658 11452
rect 19412 11398 19414 11450
rect 19594 11398 19596 11450
rect 19350 11396 19356 11398
rect 19412 11396 19436 11398
rect 19492 11396 19516 11398
rect 19572 11396 19596 11398
rect 19652 11396 19658 11398
rect 19350 11387 19658 11396
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 20456 11150 20484 13382
rect 20628 13330 20680 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20548 12986 20576 13262
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20640 12866 20668 13126
rect 20732 12986 20760 13806
rect 20824 13530 20852 13926
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21100 13530 21128 13874
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 20850 13084 21158 13093
rect 20850 13082 20856 13084
rect 20912 13082 20936 13084
rect 20992 13082 21016 13084
rect 21072 13082 21096 13084
rect 21152 13082 21158 13084
rect 20912 13030 20914 13082
rect 21094 13030 21096 13082
rect 20850 13028 20856 13030
rect 20912 13028 20936 13030
rect 20992 13028 21016 13030
rect 21072 13028 21096 13030
rect 21152 13028 21158 13030
rect 20850 13019 21158 13028
rect 21192 12986 21220 13194
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21284 12866 21312 13806
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13394 21404 13670
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21468 13274 21496 14198
rect 21560 13326 21588 14991
rect 21652 14958 21680 17682
rect 21836 17610 21864 19654
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22112 18834 22140 19110
rect 22204 18850 22232 20198
rect 22350 20156 22658 20165
rect 22350 20154 22356 20156
rect 22412 20154 22436 20156
rect 22492 20154 22516 20156
rect 22572 20154 22596 20156
rect 22652 20154 22658 20156
rect 22412 20102 22414 20154
rect 22594 20102 22596 20154
rect 22350 20100 22356 20102
rect 22412 20100 22436 20102
rect 22492 20100 22516 20102
rect 22572 20100 22596 20102
rect 22652 20100 22658 20102
rect 22350 20091 22658 20100
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22350 19068 22658 19077
rect 22350 19066 22356 19068
rect 22412 19066 22436 19068
rect 22492 19066 22516 19068
rect 22572 19066 22596 19068
rect 22652 19066 22658 19068
rect 22412 19014 22414 19066
rect 22594 19014 22596 19066
rect 22350 19012 22356 19014
rect 22412 19012 22436 19014
rect 22492 19012 22516 19014
rect 22572 19012 22596 19014
rect 22652 19012 22658 19014
rect 22350 19003 22658 19012
rect 22756 18850 22784 19722
rect 22848 18970 22876 19790
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22940 18902 22968 19246
rect 22100 18828 22152 18834
rect 22204 18822 22324 18850
rect 22100 18770 22152 18776
rect 22296 18630 22324 18822
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22572 18822 22784 18850
rect 22928 18896 22980 18902
rect 22928 18838 22980 18844
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21744 15162 21772 16594
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21836 15978 21864 16526
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21836 15094 21864 15914
rect 21928 15586 21956 15982
rect 22020 15722 22048 18090
rect 22112 17542 22140 18566
rect 22388 18193 22416 18770
rect 22374 18184 22430 18193
rect 22374 18119 22430 18128
rect 22572 18086 22600 18822
rect 22744 18760 22796 18766
rect 22664 18708 22744 18714
rect 22664 18702 22796 18708
rect 22664 18686 22784 18702
rect 22664 18426 22692 18686
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22664 18290 22692 18362
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22350 17980 22658 17989
rect 22350 17978 22356 17980
rect 22412 17978 22436 17980
rect 22492 17978 22516 17980
rect 22572 17978 22596 17980
rect 22652 17978 22658 17980
rect 22412 17926 22414 17978
rect 22594 17926 22596 17978
rect 22350 17924 22356 17926
rect 22412 17924 22436 17926
rect 22492 17924 22516 17926
rect 22572 17924 22596 17926
rect 22652 17924 22658 17926
rect 22350 17915 22658 17924
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 16794 22140 17478
rect 22296 17338 22324 17614
rect 22756 17610 22784 18566
rect 22940 18222 22968 18838
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22928 18080 22980 18086
rect 22848 18028 22928 18034
rect 22848 18022 22980 18028
rect 22848 18006 22968 18022
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22350 16892 22658 16901
rect 22350 16890 22356 16892
rect 22412 16890 22436 16892
rect 22492 16890 22516 16892
rect 22572 16890 22596 16892
rect 22652 16890 22658 16892
rect 22412 16838 22414 16890
rect 22594 16838 22596 16890
rect 22350 16836 22356 16838
rect 22412 16836 22436 16838
rect 22492 16836 22516 16838
rect 22572 16836 22596 16838
rect 22652 16836 22658 16838
rect 22350 16827 22658 16836
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22204 16182 22232 16594
rect 22192 16176 22244 16182
rect 22192 16118 22244 16124
rect 22350 15804 22658 15813
rect 22350 15802 22356 15804
rect 22412 15802 22436 15804
rect 22492 15802 22516 15804
rect 22572 15802 22596 15804
rect 22652 15802 22658 15804
rect 22412 15750 22414 15802
rect 22594 15750 22596 15802
rect 22350 15748 22356 15750
rect 22412 15748 22436 15750
rect 22492 15748 22516 15750
rect 22572 15748 22596 15750
rect 22652 15748 22658 15750
rect 22350 15739 22658 15748
rect 22020 15694 22232 15722
rect 21928 15558 22048 15586
rect 22204 15570 22232 15694
rect 22848 15638 22876 18006
rect 23032 16454 23060 19790
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23124 19446 23152 19654
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 23124 18154 23152 19246
rect 23112 18148 23164 18154
rect 23112 18090 23164 18096
rect 23124 17882 23152 18090
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23216 17270 23244 19654
rect 23308 17785 23336 20402
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23492 19242 23520 20198
rect 23676 19825 23704 20402
rect 23756 19848 23808 19854
rect 23662 19816 23718 19825
rect 23756 19790 23808 19796
rect 23662 19751 23718 19760
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23572 19168 23624 19174
rect 23570 19136 23572 19145
rect 23624 19136 23626 19145
rect 23570 19071 23626 19080
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23294 17776 23350 17785
rect 23294 17711 23350 17720
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23400 16561 23428 17478
rect 23492 17338 23520 18158
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23492 16658 23520 17274
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23386 16552 23442 16561
rect 23386 16487 23442 16496
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 23676 15910 23704 19654
rect 23768 17105 23796 19790
rect 23850 19612 24158 19621
rect 23850 19610 23856 19612
rect 23912 19610 23936 19612
rect 23992 19610 24016 19612
rect 24072 19610 24096 19612
rect 24152 19610 24158 19612
rect 23912 19558 23914 19610
rect 24094 19558 24096 19610
rect 23850 19556 23856 19558
rect 23912 19556 23936 19558
rect 23992 19556 24016 19558
rect 24072 19556 24096 19558
rect 24152 19556 24158 19558
rect 23850 19547 24158 19556
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 23850 18524 24158 18533
rect 23850 18522 23856 18524
rect 23912 18522 23936 18524
rect 23992 18522 24016 18524
rect 24072 18522 24096 18524
rect 24152 18522 24158 18524
rect 23912 18470 23914 18522
rect 24094 18470 24096 18522
rect 23850 18468 23856 18470
rect 23912 18468 23936 18470
rect 23992 18468 24016 18470
rect 24072 18468 24096 18470
rect 24152 18468 24158 18470
rect 23850 18459 24158 18468
rect 24320 18465 24348 18566
rect 24306 18456 24362 18465
rect 24306 18391 24362 18400
rect 23850 17436 24158 17445
rect 23850 17434 23856 17436
rect 23912 17434 23936 17436
rect 23992 17434 24016 17436
rect 24072 17434 24096 17436
rect 24152 17434 24158 17436
rect 23912 17382 23914 17434
rect 24094 17382 24096 17434
rect 23850 17380 23856 17382
rect 23912 17380 23936 17382
rect 23992 17380 24016 17382
rect 24072 17380 24096 17382
rect 24152 17380 24158 17382
rect 23850 17371 24158 17380
rect 23754 17096 23810 17105
rect 23754 17031 23810 17040
rect 23850 16348 24158 16357
rect 23850 16346 23856 16348
rect 23912 16346 23936 16348
rect 23992 16346 24016 16348
rect 24072 16346 24096 16348
rect 24152 16346 24158 16348
rect 23912 16294 23914 16346
rect 24094 16294 24096 16346
rect 23850 16292 23856 16294
rect 23912 16292 23936 16294
rect 23992 16292 24016 16294
rect 24072 16292 24096 16294
rect 24152 16292 24158 16294
rect 23850 16283 24158 16292
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23386 15736 23442 15745
rect 23296 15700 23348 15706
rect 23386 15671 23442 15680
rect 23296 15642 23348 15648
rect 22284 15632 22336 15638
rect 22282 15600 22284 15609
rect 22836 15632 22888 15638
rect 22336 15600 22338 15609
rect 22020 15502 22048 15558
rect 22192 15564 22244 15570
rect 22836 15574 22888 15580
rect 22282 15535 22338 15544
rect 22192 15506 22244 15512
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21652 13462 21680 14894
rect 21836 14414 21864 15030
rect 21928 14890 21956 15438
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21928 14550 21956 14826
rect 21916 14544 21968 14550
rect 21916 14486 21968 14492
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21640 13456 21692 13462
rect 21692 13404 21772 13410
rect 21640 13398 21772 13404
rect 21652 13382 21772 13398
rect 20640 12838 20760 12866
rect 20732 12442 20760 12838
rect 21192 12838 21312 12866
rect 21376 13246 21496 13274
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21640 13252 21692 13258
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 21100 12102 21128 12718
rect 21192 12714 21220 12838
rect 21272 12776 21324 12782
rect 21376 12730 21404 13246
rect 21640 13194 21692 13200
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21324 12724 21404 12730
rect 21272 12718 21404 12724
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21284 12702 21404 12718
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20850 11996 21158 12005
rect 20850 11994 20856 11996
rect 20912 11994 20936 11996
rect 20992 11994 21016 11996
rect 21072 11994 21096 11996
rect 21152 11994 21158 11996
rect 20912 11942 20914 11994
rect 21094 11942 21096 11994
rect 20850 11940 20856 11942
rect 20912 11940 20936 11942
rect 20992 11940 21016 11942
rect 21072 11940 21096 11942
rect 21152 11940 21158 11942
rect 20850 11931 21158 11940
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 17850 10908 18158 10917
rect 17850 10906 17856 10908
rect 17912 10906 17936 10908
rect 17992 10906 18016 10908
rect 18072 10906 18096 10908
rect 18152 10906 18158 10908
rect 17912 10854 17914 10906
rect 18094 10854 18096 10906
rect 17850 10852 17856 10854
rect 17912 10852 17936 10854
rect 17992 10852 18016 10854
rect 18072 10852 18096 10854
rect 18152 10852 18158 10854
rect 17850 10843 18158 10852
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 17144 8634 17172 9862
rect 17328 9722 17356 10406
rect 19350 10364 19658 10373
rect 19350 10362 19356 10364
rect 19412 10362 19436 10364
rect 19492 10362 19516 10364
rect 19572 10362 19596 10364
rect 19652 10362 19658 10364
rect 19412 10310 19414 10362
rect 19594 10310 19596 10362
rect 19350 10308 19356 10310
rect 19412 10308 19436 10310
rect 19492 10308 19516 10310
rect 19572 10308 19596 10310
rect 19652 10308 19658 10310
rect 19350 10299 19658 10308
rect 19720 10266 19748 10610
rect 19812 10470 19840 11086
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 17850 9820 18158 9829
rect 17850 9818 17856 9820
rect 17912 9818 17936 9820
rect 17992 9818 18016 9820
rect 18072 9818 18096 9820
rect 18152 9818 18158 9820
rect 17912 9766 17914 9818
rect 18094 9766 18096 9818
rect 17850 9764 17856 9766
rect 17912 9764 17936 9766
rect 17992 9764 18016 9766
rect 18072 9764 18096 9766
rect 18152 9764 18158 9766
rect 17850 9755 18158 9764
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 18524 9586 18552 10066
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 19076 9574 19656 9602
rect 19812 9586 19840 10406
rect 20088 10266 20116 11018
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20732 10062 20760 11222
rect 20850 10908 21158 10917
rect 20850 10906 20856 10908
rect 20912 10906 20936 10908
rect 20992 10906 21016 10908
rect 21072 10906 21096 10908
rect 21152 10906 21158 10908
rect 20912 10854 20914 10906
rect 21094 10854 21096 10906
rect 20850 10852 20856 10854
rect 20912 10852 20936 10854
rect 20992 10852 21016 10854
rect 21072 10852 21096 10854
rect 21152 10852 21158 10854
rect 20850 10843 21158 10852
rect 21192 10810 21220 11630
rect 21284 11558 21312 12702
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21376 12306 21404 12582
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21468 11898 21496 12786
rect 21560 12238 21588 13126
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21652 12102 21680 13194
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21284 11218 21312 11494
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20916 10198 20944 10406
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 21192 10130 21220 10746
rect 21284 10742 21312 10950
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20850 9820 21158 9829
rect 20850 9818 20856 9820
rect 20912 9818 20936 9820
rect 20992 9818 21016 9820
rect 21072 9818 21096 9820
rect 21152 9818 21158 9820
rect 20912 9766 20914 9818
rect 21094 9766 21096 9818
rect 20850 9764 20856 9766
rect 20912 9764 20936 9766
rect 20992 9764 21016 9766
rect 21072 9764 21096 9766
rect 21152 9764 21158 9766
rect 20850 9755 21158 9764
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 15198 8256 15254 8265
rect 15198 8191 15254 8200
rect 14556 7744 14608 7750
rect 14608 7704 14688 7732
rect 14556 7686 14608 7692
rect 14476 7398 14596 7426
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14476 6798 14504 7278
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14476 6390 14504 6734
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 13350 2748 13658 2757
rect 13350 2746 13356 2748
rect 13412 2746 13436 2748
rect 13492 2746 13516 2748
rect 13572 2746 13596 2748
rect 13652 2746 13658 2748
rect 14200 2746 14412 2774
rect 13412 2694 13414 2746
rect 13594 2694 13596 2746
rect 13350 2692 13356 2694
rect 13412 2692 13436 2694
rect 13492 2692 13516 2694
rect 13572 2692 13596 2694
rect 13652 2692 13658 2694
rect 13350 2683 13658 2692
rect 14384 2650 14412 2746
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14568 2446 14596 7398
rect 14660 6322 14688 7704
rect 14850 7644 15158 7653
rect 14850 7642 14856 7644
rect 14912 7642 14936 7644
rect 14992 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15158 7644
rect 14912 7590 14914 7642
rect 15094 7590 15096 7642
rect 14850 7588 14856 7590
rect 14912 7588 14936 7590
rect 14992 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15158 7590
rect 14850 7579 15158 7588
rect 15212 7478 15240 8191
rect 16350 8188 16658 8197
rect 16350 8186 16356 8188
rect 16412 8186 16436 8188
rect 16492 8186 16516 8188
rect 16572 8186 16596 8188
rect 16652 8186 16658 8188
rect 16412 8134 16414 8186
rect 16594 8134 16596 8186
rect 16350 8132 16356 8134
rect 16412 8132 16436 8134
rect 16492 8132 16516 8134
rect 16572 8132 16596 8134
rect 16652 8132 16658 8134
rect 16350 8123 16658 8132
rect 17236 8022 17264 9454
rect 18248 8906 18276 9454
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 17788 8090 17816 8842
rect 18432 8838 18460 9454
rect 19076 9450 19104 9574
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 17850 8732 18158 8741
rect 17850 8730 17856 8732
rect 17912 8730 17936 8732
rect 17992 8730 18016 8732
rect 18072 8730 18096 8732
rect 18152 8730 18158 8732
rect 17912 8678 17914 8730
rect 18094 8678 18096 8730
rect 17850 8676 17856 8678
rect 17912 8676 17936 8678
rect 17992 8676 18016 8678
rect 18072 8676 18096 8678
rect 18152 8676 18158 8678
rect 17850 8667 18158 8676
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17224 8016 17276 8022
rect 17880 7970 17908 8366
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17224 7958 17276 7964
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14850 6556 15158 6565
rect 14850 6554 14856 6556
rect 14912 6554 14936 6556
rect 14992 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15158 6556
rect 14912 6502 14914 6554
rect 15094 6502 15096 6554
rect 14850 6500 14856 6502
rect 14912 6500 14936 6502
rect 14992 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15158 6502
rect 14850 6491 15158 6500
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14660 3602 14688 6258
rect 15212 6254 15240 6666
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 14850 5468 15158 5477
rect 14850 5466 14856 5468
rect 14912 5466 14936 5468
rect 14992 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15158 5468
rect 14912 5414 14914 5466
rect 15094 5414 15096 5466
rect 14850 5412 14856 5414
rect 14912 5412 14936 5414
rect 14992 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15158 5414
rect 14850 5403 15158 5412
rect 15304 5370 15332 6598
rect 15488 6186 15516 7278
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15580 6934 15608 7210
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15488 5914 15516 6122
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5574 15516 5714
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15488 5234 15516 5510
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 14850 4380 15158 4389
rect 14850 4378 14856 4380
rect 14912 4378 14936 4380
rect 14992 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15158 4380
rect 14912 4326 14914 4378
rect 15094 4326 15096 4378
rect 14850 4324 14856 4326
rect 14912 4324 14936 4326
rect 14992 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15158 4326
rect 14850 4315 15158 4324
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14752 3505 14780 4014
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 14936 3534 14964 3878
rect 14924 3528 14976 3534
rect 14738 3496 14794 3505
rect 14924 3470 14976 3476
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 14738 3431 14794 3440
rect 14752 3194 14780 3431
rect 14850 3292 15158 3301
rect 14850 3290 14856 3292
rect 14912 3290 14936 3292
rect 14992 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15158 3292
rect 14912 3238 14914 3290
rect 15094 3238 15096 3290
rect 14850 3236 14856 3238
rect 14912 3236 14936 3238
rect 14992 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15158 3238
rect 14850 3227 15158 3236
rect 15212 3194 15240 3470
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15304 3126 15332 3470
rect 15396 3194 15424 3878
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15304 2650 15332 3062
rect 15580 2990 15608 6870
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 4690 15700 6802
rect 15764 6458 15792 7142
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 16040 6390 16068 6598
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4146 15700 4626
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3058 15792 3878
rect 15948 3534 15976 4082
rect 16040 3738 16068 6054
rect 16132 5234 16160 7142
rect 16350 7100 16658 7109
rect 16350 7098 16356 7100
rect 16412 7098 16436 7100
rect 16492 7098 16516 7100
rect 16572 7098 16596 7100
rect 16652 7098 16658 7100
rect 16412 7046 16414 7098
rect 16594 7046 16596 7098
rect 16350 7044 16356 7046
rect 16412 7044 16436 7046
rect 16492 7044 16516 7046
rect 16572 7044 16596 7046
rect 16652 7044 16658 7046
rect 16350 7035 16658 7044
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16224 5370 16252 6598
rect 16350 6012 16658 6021
rect 16350 6010 16356 6012
rect 16412 6010 16436 6012
rect 16492 6010 16516 6012
rect 16572 6010 16596 6012
rect 16652 6010 16658 6012
rect 16412 5958 16414 6010
rect 16594 5958 16596 6010
rect 16350 5956 16356 5958
rect 16412 5956 16436 5958
rect 16492 5956 16516 5958
rect 16572 5956 16596 5958
rect 16652 5956 16658 5958
rect 16350 5947 16658 5956
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16316 5012 16344 5646
rect 16776 5370 16804 6734
rect 16868 6186 16896 7346
rect 17236 7342 17264 7958
rect 17788 7942 17908 7970
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16868 5250 16896 6122
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5846 16988 6054
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16776 5234 16896 5250
rect 16764 5228 16896 5234
rect 16816 5222 16896 5228
rect 16764 5170 16816 5176
rect 16224 4984 16344 5012
rect 16224 4214 16252 4984
rect 16350 4924 16658 4933
rect 16350 4922 16356 4924
rect 16412 4922 16436 4924
rect 16492 4922 16516 4924
rect 16572 4922 16596 4924
rect 16652 4922 16658 4924
rect 16412 4870 16414 4922
rect 16594 4870 16596 4922
rect 16350 4868 16356 4870
rect 16412 4868 16436 4870
rect 16492 4868 16516 4870
rect 16572 4868 16596 4870
rect 16652 4868 16658 4870
rect 16350 4859 16658 4868
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16132 3602 16160 3946
rect 16350 3836 16658 3845
rect 16350 3834 16356 3836
rect 16412 3834 16436 3836
rect 16492 3834 16516 3836
rect 16572 3834 16596 3836
rect 16652 3834 16658 3836
rect 16412 3782 16414 3834
rect 16594 3782 16596 3834
rect 16350 3780 16356 3782
rect 16412 3780 16436 3782
rect 16492 3780 16516 3782
rect 16572 3780 16596 3782
rect 16652 3780 16658 3782
rect 16350 3771 16658 3780
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15936 3528 15988 3534
rect 16212 3528 16264 3534
rect 15936 3470 15988 3476
rect 16210 3496 16212 3505
rect 16264 3496 16266 3505
rect 16210 3431 16266 3440
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16350 2748 16658 2757
rect 16350 2746 16356 2748
rect 16412 2746 16436 2748
rect 16492 2746 16516 2748
rect 16572 2746 16596 2748
rect 16652 2746 16658 2748
rect 16412 2694 16414 2746
rect 16594 2694 16596 2746
rect 16350 2692 16356 2694
rect 16412 2692 16436 2694
rect 16492 2692 16516 2694
rect 16572 2692 16596 2694
rect 16652 2692 16658 2694
rect 16350 2683 16658 2692
rect 16776 2650 16804 5170
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16868 4010 16896 4490
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16960 3194 16988 4490
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17052 3602 17080 4422
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17144 3482 17172 4082
rect 17052 3454 17172 3482
rect 17052 3194 17080 3454
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17052 3058 17080 3130
rect 17144 3058 17172 3334
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17236 2990 17264 7278
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17512 5370 17540 6598
rect 17604 6458 17632 6734
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17604 5710 17632 6394
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17696 5574 17724 7346
rect 17788 7274 17816 7942
rect 17972 7886 18000 8230
rect 18064 7954 18092 8502
rect 18432 7954 18460 8774
rect 18892 8634 18920 9318
rect 19076 9110 19104 9386
rect 19168 9178 19196 9386
rect 19260 9178 19288 9454
rect 19628 9450 19656 9574
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19350 9276 19658 9285
rect 19350 9274 19356 9276
rect 19412 9274 19436 9276
rect 19492 9274 19516 9276
rect 19572 9274 19596 9276
rect 19652 9274 19658 9276
rect 19412 9222 19414 9274
rect 19594 9222 19596 9274
rect 19350 9220 19356 9222
rect 19412 9220 19436 9222
rect 19492 9220 19516 9222
rect 19572 9220 19596 9222
rect 19652 9220 19658 9222
rect 19350 9211 19658 9220
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19812 8974 19840 9522
rect 21284 9450 21312 10202
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21376 9466 21404 9998
rect 21468 9586 21496 11222
rect 21652 10810 21680 11494
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21744 10606 21772 13382
rect 21836 13326 21864 14350
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21836 12918 21864 13262
rect 21928 13190 21956 13806
rect 22100 13728 22152 13734
rect 22098 13696 22100 13705
rect 22152 13696 22154 13705
rect 22098 13631 22154 13640
rect 22204 13546 22232 15506
rect 22350 14716 22658 14725
rect 22350 14714 22356 14716
rect 22412 14714 22436 14716
rect 22492 14714 22516 14716
rect 22572 14714 22596 14716
rect 22652 14714 22658 14716
rect 22412 14662 22414 14714
rect 22594 14662 22596 14714
rect 22350 14660 22356 14662
rect 22412 14660 22436 14662
rect 22492 14660 22516 14662
rect 22572 14660 22596 14662
rect 22652 14660 22658 14662
rect 22350 14651 22658 14660
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22480 14074 22508 14350
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22848 13954 22876 15574
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22940 14074 22968 14962
rect 23032 14822 23060 15438
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 22848 13926 22968 13954
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22350 13628 22658 13637
rect 22350 13626 22356 13628
rect 22412 13626 22436 13628
rect 22492 13626 22516 13628
rect 22572 13626 22596 13628
rect 22652 13626 22658 13628
rect 22412 13574 22414 13626
rect 22594 13574 22596 13626
rect 22350 13572 22356 13574
rect 22412 13572 22436 13574
rect 22492 13572 22516 13574
rect 22572 13572 22596 13574
rect 22652 13572 22658 13574
rect 22350 13563 22658 13572
rect 22204 13518 22324 13546
rect 22296 13274 22324 13518
rect 22192 13252 22244 13258
rect 22296 13246 22508 13274
rect 22192 13194 22244 13200
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21824 12912 21876 12918
rect 21824 12854 21876 12860
rect 21836 12306 21864 12854
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21836 10130 21864 11290
rect 21928 10674 21956 12582
rect 22112 12238 22140 12582
rect 22204 12442 22232 13194
rect 22480 12850 22508 13246
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22756 12850 22784 13126
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22350 12540 22658 12549
rect 22350 12538 22356 12540
rect 22412 12538 22436 12540
rect 22492 12538 22516 12540
rect 22572 12538 22596 12540
rect 22652 12538 22658 12540
rect 22412 12486 22414 12538
rect 22594 12486 22596 12538
rect 22350 12484 22356 12486
rect 22412 12484 22436 12486
rect 22492 12484 22516 12486
rect 22572 12484 22596 12486
rect 22652 12484 22658 12486
rect 22350 12475 22658 12484
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22848 12170 22876 13670
rect 22940 12782 22968 13926
rect 23032 13870 23060 14758
rect 23124 14618 23152 15438
rect 23308 15026 23336 15642
rect 23400 15162 23428 15671
rect 23850 15260 24158 15269
rect 23850 15258 23856 15260
rect 23912 15258 23936 15260
rect 23992 15258 24016 15260
rect 24072 15258 24096 15260
rect 24152 15258 24158 15260
rect 23912 15206 23914 15258
rect 24094 15206 24096 15258
rect 23850 15204 23856 15206
rect 23912 15204 23936 15206
rect 23992 15204 24016 15206
rect 24072 15204 24096 15206
rect 24152 15204 24158 15206
rect 23850 15195 24158 15204
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23570 14376 23626 14385
rect 23570 14311 23626 14320
rect 23584 14278 23612 14311
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23850 14172 24158 14181
rect 23850 14170 23856 14172
rect 23912 14170 23936 14172
rect 23992 14170 24016 14172
rect 24072 14170 24096 14172
rect 24152 14170 24158 14172
rect 23912 14118 23914 14170
rect 24094 14118 24096 14170
rect 23850 14116 23856 14118
rect 23912 14116 23936 14118
rect 23992 14116 24016 14118
rect 24072 14116 24096 14118
rect 24152 14116 24158 14118
rect 23850 14107 24158 14116
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23662 13696 23718 13705
rect 23662 13631 23718 13640
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 23216 12238 23244 12922
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23308 12442 23336 12786
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11762 22232 12038
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22848 11694 22876 12106
rect 23308 11762 23336 12378
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22350 11452 22658 11461
rect 22350 11450 22356 11452
rect 22412 11450 22436 11452
rect 22492 11450 22516 11452
rect 22572 11450 22596 11452
rect 22652 11450 22658 11452
rect 22412 11398 22414 11450
rect 22594 11398 22596 11450
rect 22350 11396 22356 11398
rect 22412 11396 22436 11398
rect 22492 11396 22516 11398
rect 22572 11396 22596 11398
rect 22652 11396 22658 11398
rect 22350 11387 22658 11396
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10742 22048 11086
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 22020 9586 22048 10678
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21548 9512 21600 9518
rect 20444 9444 20496 9450
rect 20444 9386 20496 9392
rect 21272 9444 21324 9450
rect 21376 9438 21496 9466
rect 21548 9454 21600 9460
rect 21272 9386 21324 9392
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19536 8634 19564 8842
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19812 8566 19840 8910
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 8090 19288 8434
rect 19904 8430 19932 8774
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19350 8188 19658 8197
rect 19350 8186 19356 8188
rect 19412 8186 19436 8188
rect 19492 8186 19516 8188
rect 19572 8186 19596 8188
rect 19652 8186 19658 8188
rect 19412 8134 19414 8186
rect 19594 8134 19596 8186
rect 19350 8132 19356 8134
rect 19412 8132 19436 8134
rect 19492 8132 19516 8134
rect 19572 8132 19596 8134
rect 19652 8132 19658 8134
rect 19350 8123 19658 8132
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19720 7954 19748 8230
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19904 7886 19932 8366
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 17850 7644 18158 7653
rect 17850 7642 17856 7644
rect 17912 7642 17936 7644
rect 17992 7642 18016 7644
rect 18072 7642 18096 7644
rect 18152 7642 18158 7644
rect 17912 7590 17914 7642
rect 18094 7590 18096 7642
rect 17850 7588 17856 7590
rect 17912 7588 17936 7590
rect 17992 7588 18016 7590
rect 18072 7588 18096 7590
rect 18152 7588 18158 7590
rect 17850 7579 18158 7588
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17972 6730 18000 7278
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 17850 6556 18158 6565
rect 17850 6554 17856 6556
rect 17912 6554 17936 6556
rect 17992 6554 18016 6556
rect 18072 6554 18096 6556
rect 18152 6554 18158 6556
rect 17912 6502 17914 6554
rect 18094 6502 18096 6554
rect 17850 6500 17856 6502
rect 17912 6500 17936 6502
rect 17992 6500 18016 6502
rect 18072 6500 18096 6502
rect 18152 6500 18158 6502
rect 17850 6491 18158 6500
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17328 4078 17356 5102
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17512 4282 17540 4966
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 17328 3126 17356 3402
rect 17420 3194 17448 4082
rect 17788 4078 17816 6054
rect 18156 5658 18184 6258
rect 18248 5778 18276 6666
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18340 5710 18368 6598
rect 18328 5704 18380 5710
rect 18156 5630 18276 5658
rect 18328 5646 18380 5652
rect 17850 5468 18158 5477
rect 17850 5466 17856 5468
rect 17912 5466 17936 5468
rect 17992 5466 18016 5468
rect 18072 5466 18096 5468
rect 18152 5466 18158 5468
rect 17912 5414 17914 5466
rect 18094 5414 18096 5466
rect 17850 5412 17856 5414
rect 17912 5412 17936 5414
rect 17992 5412 18016 5414
rect 18072 5412 18096 5414
rect 18152 5412 18158 5414
rect 17850 5403 18158 5412
rect 18248 5250 18276 5630
rect 18248 5222 18368 5250
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 17850 4380 18158 4389
rect 17850 4378 17856 4380
rect 17912 4378 17936 4380
rect 17992 4378 18016 4380
rect 18072 4378 18096 4380
rect 18152 4378 18158 4380
rect 17912 4326 17914 4378
rect 18094 4326 18096 4378
rect 17850 4324 17856 4326
rect 17912 4324 17936 4326
rect 17992 4324 18016 4326
rect 18072 4324 18096 4326
rect 18152 4324 18158 4326
rect 17850 4315 18158 4324
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17788 3534 17816 4014
rect 18248 3738 18276 5102
rect 18340 4690 18368 5222
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17788 3058 17816 3470
rect 17850 3292 18158 3301
rect 17850 3290 17856 3292
rect 17912 3290 17936 3292
rect 17992 3290 18016 3292
rect 18072 3290 18096 3292
rect 18152 3290 18158 3292
rect 17912 3238 17914 3290
rect 18094 3238 18096 3290
rect 17850 3236 17856 3238
rect 17912 3236 17936 3238
rect 17992 3236 18016 3238
rect 18072 3236 18096 3238
rect 18152 3236 18158 3238
rect 17850 3227 18158 3236
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17512 2514 17540 2790
rect 18340 2650 18368 4082
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 2850 2204 3158 2213
rect 2850 2202 2856 2204
rect 2912 2202 2936 2204
rect 2992 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3158 2204
rect 2912 2150 2914 2202
rect 3094 2150 3096 2202
rect 2850 2148 2856 2150
rect 2912 2148 2936 2150
rect 2992 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3158 2150
rect 2850 2139 3158 2148
rect 5736 1306 5764 2382
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5850 2204 6158 2213
rect 5850 2202 5856 2204
rect 5912 2202 5936 2204
rect 5992 2202 6016 2204
rect 6072 2202 6096 2204
rect 6152 2202 6158 2204
rect 5912 2150 5914 2202
rect 6094 2150 6096 2202
rect 5850 2148 5856 2150
rect 5912 2148 5936 2150
rect 5992 2148 6016 2150
rect 6072 2148 6096 2150
rect 6152 2148 6158 2150
rect 5850 2139 6158 2148
rect 5736 1278 5856 1306
rect 5828 400 5856 1278
rect 6472 400 6500 2246
rect 7116 400 7144 2314
rect 7760 400 7788 2314
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 400 8432 2246
rect 8850 2204 9158 2213
rect 8850 2202 8856 2204
rect 8912 2202 8936 2204
rect 8992 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9158 2204
rect 8912 2150 8914 2202
rect 9094 2150 9096 2202
rect 8850 2148 8856 2150
rect 8912 2148 8936 2150
rect 8992 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9158 2150
rect 8850 2139 9158 2148
rect 9232 1306 9260 2382
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9048 1278 9260 1306
rect 9048 400 9076 1278
rect 9692 400 9720 2314
rect 10336 400 10364 2382
rect 11624 400 11652 2382
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 11850 2204 12158 2213
rect 11850 2202 11856 2204
rect 11912 2202 11936 2204
rect 11992 2202 12016 2204
rect 12072 2202 12096 2204
rect 12152 2202 12158 2204
rect 11912 2150 11914 2202
rect 12094 2150 12096 2202
rect 11850 2148 11856 2150
rect 11912 2148 11936 2150
rect 11992 2148 12016 2150
rect 12072 2148 12096 2150
rect 12152 2148 12158 2150
rect 11850 2139 12158 2148
rect 12268 400 12296 2314
rect 14200 400 14228 2382
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 1170 14780 2246
rect 14850 2204 15158 2213
rect 14850 2202 14856 2204
rect 14912 2202 14936 2204
rect 14992 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15158 2204
rect 14912 2150 14914 2202
rect 15094 2150 15096 2202
rect 14850 2148 14856 2150
rect 14912 2148 14936 2150
rect 14992 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15158 2150
rect 14850 2139 15158 2148
rect 14752 1142 14872 1170
rect 14844 400 14872 1142
rect 15488 400 15516 2382
rect 16132 400 16160 2382
rect 18432 2378 18460 7142
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18524 5914 18552 6258
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18800 5710 18828 7142
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18892 6390 18920 6802
rect 19076 6730 19104 7346
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19350 7100 19658 7109
rect 19350 7098 19356 7100
rect 19412 7098 19436 7100
rect 19492 7098 19516 7100
rect 19572 7098 19596 7100
rect 19652 7098 19658 7100
rect 19412 7046 19414 7098
rect 19594 7046 19596 7098
rect 19350 7044 19356 7046
rect 19412 7044 19436 7046
rect 19492 7044 19516 7046
rect 19572 7044 19596 7046
rect 19652 7044 19658 7046
rect 19350 7035 19658 7044
rect 19720 6866 19748 7142
rect 19812 6866 19840 7482
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 5914 19012 6258
rect 19720 6254 19748 6666
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19350 6012 19658 6021
rect 19350 6010 19356 6012
rect 19412 6010 19436 6012
rect 19492 6010 19516 6012
rect 19572 6010 19596 6012
rect 19652 6010 19658 6012
rect 19412 5958 19414 6010
rect 19594 5958 19596 6010
rect 19350 5956 19356 5958
rect 19412 5956 19436 5958
rect 19492 5956 19516 5958
rect 19572 5956 19596 5958
rect 19652 5956 19658 5958
rect 19350 5947 19658 5956
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 19720 5778 19748 6190
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19350 4924 19658 4933
rect 19350 4922 19356 4924
rect 19412 4922 19436 4924
rect 19492 4922 19516 4924
rect 19572 4922 19596 4924
rect 19652 4922 19658 4924
rect 19412 4870 19414 4922
rect 19594 4870 19596 4922
rect 19350 4868 19356 4870
rect 19412 4868 19436 4870
rect 19492 4868 19516 4870
rect 19572 4868 19596 4870
rect 19652 4868 19658 4870
rect 19350 4859 19658 4868
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 18892 3534 18920 4422
rect 19536 4078 19564 4422
rect 19720 4146 19748 5034
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19350 3836 19658 3845
rect 19350 3834 19356 3836
rect 19412 3834 19436 3836
rect 19492 3834 19516 3836
rect 19572 3834 19596 3836
rect 19652 3834 19658 3836
rect 19412 3782 19414 3834
rect 19594 3782 19596 3834
rect 19350 3780 19356 3782
rect 19412 3780 19436 3782
rect 19492 3780 19516 3782
rect 19572 3780 19596 3782
rect 19652 3780 19658 3782
rect 19350 3771 19658 3780
rect 19720 3738 19748 4082
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 18708 3126 18736 3334
rect 19720 3194 19748 3334
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19812 3126 19840 4626
rect 19904 4010 19932 5850
rect 19996 5302 20024 7890
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20088 6934 20116 7278
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20088 6458 20116 6870
rect 20456 6866 20484 9386
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20732 8498 20760 9114
rect 21192 8974 21220 9318
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21468 8906 21496 9438
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 20850 8732 21158 8741
rect 20850 8730 20856 8732
rect 20912 8730 20936 8732
rect 20992 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21158 8732
rect 20912 8678 20914 8730
rect 21094 8678 21096 8730
rect 20850 8676 20856 8678
rect 20912 8676 20936 8678
rect 20992 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21158 8678
rect 20850 8667 21158 8676
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20640 8401 20668 8434
rect 20626 8392 20682 8401
rect 20626 8327 20682 8336
rect 20720 8356 20772 8362
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20548 7546 20576 7890
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 6882 20668 8327
rect 20720 8298 20772 8304
rect 20732 8090 20760 8298
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 21088 7744 21140 7750
rect 21140 7704 21220 7732
rect 21088 7686 21140 7692
rect 20732 7546 20760 7686
rect 20850 7644 21158 7653
rect 20850 7642 20856 7644
rect 20912 7642 20936 7644
rect 20992 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21158 7644
rect 20912 7590 20914 7642
rect 21094 7590 21096 7642
rect 20850 7588 20856 7590
rect 20912 7588 20936 7590
rect 20992 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21158 7590
rect 20850 7579 21158 7588
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20732 7392 20760 7482
rect 20812 7404 20864 7410
rect 20732 7364 20812 7392
rect 20812 7346 20864 7352
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20444 6860 20496 6866
rect 20640 6854 20760 6882
rect 20916 6866 20944 6938
rect 20444 6802 20496 6808
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20180 6390 20208 6734
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20456 5846 20484 6802
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20732 5710 20760 6854
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20850 6556 21158 6565
rect 20850 6554 20856 6556
rect 20912 6554 20936 6556
rect 20992 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21158 6556
rect 20912 6502 20914 6554
rect 21094 6502 21096 6554
rect 20850 6500 20856 6502
rect 20912 6500 20936 6502
rect 20992 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21158 6502
rect 20850 6491 21158 6500
rect 21192 6322 21220 7704
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21284 5914 21312 7822
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21376 6458 21404 7346
rect 21468 6934 21496 8842
rect 21560 8090 21588 9454
rect 22020 9110 22048 9522
rect 22112 9382 22140 10610
rect 22350 10364 22658 10373
rect 22350 10362 22356 10364
rect 22412 10362 22436 10364
rect 22492 10362 22516 10364
rect 22572 10362 22596 10364
rect 22652 10362 22658 10364
rect 22412 10310 22414 10362
rect 22594 10310 22596 10362
rect 22350 10308 22356 10310
rect 22412 10308 22436 10310
rect 22492 10308 22516 10310
rect 22572 10308 22596 10310
rect 22652 10308 22658 10310
rect 22350 10299 22658 10308
rect 23032 10266 23060 10950
rect 23400 10810 23428 13262
rect 23492 12782 23520 13466
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23572 12368 23624 12374
rect 23570 12336 23572 12345
rect 23624 12336 23626 12345
rect 23570 12271 23626 12280
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23492 11665 23520 11766
rect 23676 11762 23704 13631
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 23850 13084 24158 13093
rect 23850 13082 23856 13084
rect 23912 13082 23936 13084
rect 23992 13082 24016 13084
rect 24072 13082 24096 13084
rect 24152 13082 24158 13084
rect 23912 13030 23914 13082
rect 24094 13030 24096 13082
rect 23850 13028 23856 13030
rect 23912 13028 23936 13030
rect 23992 13028 24016 13030
rect 24072 13028 24096 13030
rect 24152 13028 24158 13030
rect 23850 13019 24158 13028
rect 24320 13025 24348 13126
rect 24306 13016 24362 13025
rect 24306 12951 24362 12960
rect 23850 11996 24158 12005
rect 23850 11994 23856 11996
rect 23912 11994 23936 11996
rect 23992 11994 24016 11996
rect 24072 11994 24096 11996
rect 24152 11994 24158 11996
rect 23912 11942 23914 11994
rect 24094 11942 24096 11994
rect 23850 11940 23856 11942
rect 23912 11940 23936 11942
rect 23992 11940 24016 11942
rect 24072 11940 24096 11942
rect 24152 11940 24158 11942
rect 23850 11931 24158 11940
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23478 11656 23534 11665
rect 23478 11591 23534 11600
rect 23850 10908 24158 10917
rect 23850 10906 23856 10908
rect 23912 10906 23936 10908
rect 23992 10906 24016 10908
rect 24072 10906 24096 10908
rect 24152 10906 24158 10908
rect 23912 10854 23914 10906
rect 24094 10854 24096 10906
rect 23850 10852 23856 10854
rect 23912 10852 23936 10854
rect 23992 10852 24016 10854
rect 24072 10852 24096 10854
rect 24152 10852 24158 10854
rect 23850 10843 24158 10852
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23294 10704 23350 10713
rect 23294 10639 23350 10648
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22204 9450 22232 9998
rect 22664 9722 22692 9998
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22204 9178 22232 9386
rect 22350 9276 22658 9285
rect 22350 9274 22356 9276
rect 22412 9274 22436 9276
rect 22492 9274 22516 9276
rect 22572 9274 22596 9276
rect 22652 9274 22658 9276
rect 22412 9222 22414 9274
rect 22594 9222 22596 9274
rect 22350 9220 22356 9222
rect 22412 9220 22436 9222
rect 22492 9220 22516 9222
rect 22572 9220 22596 9222
rect 22652 9220 22658 9222
rect 22350 9211 22658 9220
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22756 8974 22784 9862
rect 22848 9625 22876 9862
rect 22834 9616 22890 9625
rect 22834 9551 22890 9560
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 22940 9178 22968 9522
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23308 9042 23336 10639
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23386 10296 23442 10305
rect 23386 10231 23442 10240
rect 23400 9450 23428 10231
rect 23584 10130 23612 10406
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23850 9820 24158 9829
rect 23850 9818 23856 9820
rect 23912 9818 23936 9820
rect 23992 9818 24016 9820
rect 24072 9818 24096 9820
rect 24152 9818 24158 9820
rect 23912 9766 23914 9818
rect 24094 9766 24096 9818
rect 23850 9764 23856 9766
rect 23912 9764 23936 9766
rect 23992 9764 24016 9766
rect 24072 9764 24096 9766
rect 24152 9764 24158 9766
rect 23850 9755 24158 9764
rect 23388 9444 23440 9450
rect 23388 9386 23440 9392
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 22744 8968 22796 8974
rect 23388 8968 23440 8974
rect 22744 8910 22796 8916
rect 23386 8936 23388 8945
rect 23440 8936 23442 8945
rect 23386 8871 23442 8880
rect 23850 8732 24158 8741
rect 23850 8730 23856 8732
rect 23912 8730 23936 8732
rect 23992 8730 24016 8732
rect 24072 8730 24096 8732
rect 24152 8730 24158 8732
rect 23912 8678 23914 8730
rect 24094 8678 24096 8730
rect 23850 8676 23856 8678
rect 23912 8676 23936 8678
rect 23992 8676 24016 8678
rect 24072 8676 24096 8678
rect 24152 8676 24158 8678
rect 23850 8667 24158 8676
rect 22350 8188 22658 8197
rect 22350 8186 22356 8188
rect 22412 8186 22436 8188
rect 22492 8186 22516 8188
rect 22572 8186 22596 8188
rect 22652 8186 22658 8188
rect 22412 8134 22414 8186
rect 22594 8134 22596 8186
rect 22350 8132 22356 8134
rect 22412 8132 22436 8134
rect 22492 8132 22516 8134
rect 22572 8132 22596 8134
rect 22652 8132 22658 8134
rect 22350 8123 22658 8132
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20088 4690 20116 5170
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19260 2446 19288 2790
rect 19812 2774 19840 3062
rect 19996 2922 20024 4558
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 20088 3942 20116 4422
rect 20272 4146 20300 4558
rect 20352 4276 20404 4282
rect 20352 4218 20404 4224
rect 20364 4146 20392 4218
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20364 3754 20392 4082
rect 20364 3738 20484 3754
rect 20364 3732 20496 3738
rect 20364 3726 20444 3732
rect 20444 3674 20496 3680
rect 20640 3058 20668 5578
rect 21468 5574 21496 6870
rect 21560 6254 21588 7482
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21652 6798 21680 7278
rect 21744 7002 21772 7278
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6322 21680 6598
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21560 5710 21588 6190
rect 21744 6186 21772 6938
rect 21836 6798 21864 7958
rect 23850 7644 24158 7653
rect 23850 7642 23856 7644
rect 23912 7642 23936 7644
rect 23992 7642 24016 7644
rect 24072 7642 24096 7644
rect 24152 7642 24158 7644
rect 23912 7590 23914 7642
rect 24094 7590 24096 7642
rect 23850 7588 23856 7590
rect 23912 7588 23936 7590
rect 23992 7588 24016 7590
rect 24072 7588 24096 7590
rect 24152 7588 24158 7590
rect 23850 7579 24158 7588
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22350 7100 22658 7109
rect 22350 7098 22356 7100
rect 22412 7098 22436 7100
rect 22492 7098 22516 7100
rect 22572 7098 22596 7100
rect 22652 7098 22658 7100
rect 22412 7046 22414 7098
rect 22594 7046 22596 7098
rect 22350 7044 22356 7046
rect 22412 7044 22436 7046
rect 22492 7044 22516 7046
rect 22572 7044 22596 7046
rect 22652 7044 22658 7046
rect 22350 7035 22658 7044
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 22848 6458 22876 7346
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23400 6905 23428 7142
rect 23386 6896 23442 6905
rect 23386 6831 23442 6840
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 23124 6390 23152 6598
rect 23850 6556 24158 6565
rect 23850 6554 23856 6556
rect 23912 6554 23936 6556
rect 23992 6554 24016 6556
rect 24072 6554 24096 6556
rect 24152 6554 24158 6556
rect 23912 6502 23914 6554
rect 24094 6502 24096 6554
rect 23850 6500 23856 6502
rect 23912 6500 23936 6502
rect 23992 6500 24016 6502
rect 24072 6500 24096 6502
rect 24152 6500 24158 6502
rect 23850 6491 24158 6500
rect 23112 6384 23164 6390
rect 23112 6326 23164 6332
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 6225 23704 6258
rect 23662 6216 23718 6225
rect 21732 6180 21784 6186
rect 23662 6151 23718 6160
rect 21732 6122 21784 6128
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22204 5846 22232 6054
rect 22350 6012 22658 6021
rect 22350 6010 22356 6012
rect 22412 6010 22436 6012
rect 22492 6010 22516 6012
rect 22572 6010 22596 6012
rect 22652 6010 22658 6012
rect 22412 5958 22414 6010
rect 22594 5958 22596 6010
rect 22350 5956 22356 5958
rect 22412 5956 22436 5958
rect 22492 5956 22516 5958
rect 22572 5956 22596 5958
rect 22652 5956 22658 5958
rect 22350 5947 22658 5956
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 20732 4078 20760 5510
rect 20850 5468 21158 5477
rect 20850 5466 20856 5468
rect 20912 5466 20936 5468
rect 20992 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21158 5468
rect 20912 5414 20914 5466
rect 21094 5414 21096 5466
rect 20850 5412 20856 5414
rect 20912 5412 20936 5414
rect 20992 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21158 5414
rect 20850 5403 21158 5412
rect 23850 5468 24158 5477
rect 23850 5466 23856 5468
rect 23912 5466 23936 5468
rect 23992 5466 24016 5468
rect 24072 5466 24096 5468
rect 24152 5466 24158 5468
rect 23912 5414 23914 5466
rect 24094 5414 24096 5466
rect 23850 5412 23856 5414
rect 23912 5412 23936 5414
rect 23992 5412 24016 5414
rect 24072 5412 24096 5414
rect 24152 5412 24158 5414
rect 23850 5403 24158 5412
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 20850 4380 21158 4389
rect 20850 4378 20856 4380
rect 20912 4378 20936 4380
rect 20992 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21158 4380
rect 20912 4326 20914 4378
rect 21094 4326 21096 4378
rect 20850 4324 20856 4326
rect 20912 4324 20936 4326
rect 20992 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21158 4326
rect 20850 4315 21158 4324
rect 21284 4282 21312 4490
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 21376 3534 21404 4558
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20850 3292 21158 3301
rect 20850 3290 20856 3292
rect 20912 3290 20936 3292
rect 20992 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21158 3292
rect 20912 3238 20914 3290
rect 21094 3238 21096 3290
rect 20850 3236 20856 3238
rect 20912 3236 20936 3238
rect 20992 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21158 3238
rect 20850 3227 21158 3236
rect 21468 3194 21496 4082
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21652 3602 21680 3878
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 21744 3534 21772 4966
rect 22350 4924 22658 4933
rect 22350 4922 22356 4924
rect 22412 4922 22436 4924
rect 22492 4922 22516 4924
rect 22572 4922 22596 4924
rect 22652 4922 22658 4924
rect 22412 4870 22414 4922
rect 22594 4870 22596 4922
rect 22350 4868 22356 4870
rect 22412 4868 22436 4870
rect 22492 4868 22516 4870
rect 22572 4868 22596 4870
rect 22652 4868 22658 4870
rect 22350 4859 22658 4868
rect 23850 4380 24158 4389
rect 23850 4378 23856 4380
rect 23912 4378 23936 4380
rect 23992 4378 24016 4380
rect 24072 4378 24096 4380
rect 24152 4378 24158 4380
rect 23912 4326 23914 4378
rect 24094 4326 24096 4378
rect 23850 4324 23856 4326
rect 23912 4324 23936 4326
rect 23992 4324 24016 4326
rect 24072 4324 24096 4326
rect 24152 4324 24158 4326
rect 23850 4315 24158 4324
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21836 3126 21864 3878
rect 22350 3836 22658 3845
rect 22350 3834 22356 3836
rect 22412 3834 22436 3836
rect 22492 3834 22516 3836
rect 22572 3834 22596 3836
rect 22652 3834 22658 3836
rect 22412 3782 22414 3834
rect 22594 3782 22596 3834
rect 22350 3780 22356 3782
rect 22412 3780 22436 3782
rect 22492 3780 22516 3782
rect 22572 3780 22596 3782
rect 22652 3780 22658 3782
rect 22350 3771 22658 3780
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19350 2748 19658 2757
rect 19350 2746 19356 2748
rect 19412 2746 19436 2748
rect 19492 2746 19516 2748
rect 19572 2746 19596 2748
rect 19652 2746 19658 2748
rect 19412 2694 19414 2746
rect 19594 2694 19596 2746
rect 19350 2692 19356 2694
rect 19412 2692 19436 2694
rect 19492 2692 19516 2694
rect 19572 2692 19596 2694
rect 19652 2692 19658 2694
rect 19350 2683 19658 2692
rect 19720 2746 19840 2774
rect 19720 2650 19748 2746
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 21928 2446 21956 3334
rect 23850 3292 24158 3301
rect 23850 3290 23856 3292
rect 23912 3290 23936 3292
rect 23992 3290 24016 3292
rect 24072 3290 24096 3292
rect 24152 3290 24158 3292
rect 23912 3238 23914 3290
rect 24094 3238 24096 3290
rect 23850 3236 23856 3238
rect 23912 3236 23936 3238
rect 23992 3236 24016 3238
rect 24072 3236 24096 3238
rect 24152 3236 24158 3238
rect 23850 3227 24158 3236
rect 22350 2748 22658 2757
rect 22350 2746 22356 2748
rect 22412 2746 22436 2748
rect 22492 2746 22516 2748
rect 22572 2746 22596 2748
rect 22652 2746 22658 2748
rect 22412 2694 22414 2746
rect 22594 2694 22596 2746
rect 22350 2692 22356 2694
rect 22412 2692 22436 2694
rect 22492 2692 22516 2694
rect 22572 2692 22596 2694
rect 22652 2692 22658 2694
rect 22350 2683 22658 2692
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 16776 400 16804 2314
rect 17420 400 17448 2314
rect 17850 2204 18158 2213
rect 17850 2202 17856 2204
rect 17912 2202 17936 2204
rect 17992 2202 18016 2204
rect 18072 2202 18096 2204
rect 18152 2202 18158 2204
rect 17912 2150 17914 2202
rect 18094 2150 18096 2202
rect 17850 2148 17856 2150
rect 17912 2148 17936 2150
rect 17992 2148 18016 2150
rect 18072 2148 18096 2150
rect 18152 2148 18158 2150
rect 17850 2139 18158 2148
rect 19352 400 19380 2382
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 20850 2204 21158 2213
rect 20850 2202 20856 2204
rect 20912 2202 20936 2204
rect 20992 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21158 2204
rect 20912 2150 20914 2202
rect 21094 2150 21096 2202
rect 20850 2148 20856 2150
rect 20912 2148 20936 2150
rect 20992 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21158 2150
rect 20850 2139 21158 2148
rect 21284 400 21312 2246
rect 23850 2204 24158 2213
rect 23850 2202 23856 2204
rect 23912 2202 23936 2204
rect 23992 2202 24016 2204
rect 24072 2202 24096 2204
rect 24152 2202 24158 2204
rect 23912 2150 23914 2202
rect 24094 2150 24096 2202
rect 23850 2148 23856 2150
rect 23912 2148 23936 2150
rect 23992 2148 24016 2150
rect 24072 2148 24096 2150
rect 24152 2148 24158 2150
rect 23850 2139 24158 2148
rect 5814 0 5870 400
rect 6458 0 6514 400
rect 7102 0 7158 400
rect 7746 0 7802 400
rect 8390 0 8446 400
rect 9034 0 9090 400
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 19338 0 19394 400
rect 21270 0 21326 400
<< via2 >>
rect 2856 25050 2912 25052
rect 2936 25050 2992 25052
rect 3016 25050 3072 25052
rect 3096 25050 3152 25052
rect 2856 24998 2902 25050
rect 2902 24998 2912 25050
rect 2936 24998 2966 25050
rect 2966 24998 2978 25050
rect 2978 24998 2992 25050
rect 3016 24998 3030 25050
rect 3030 24998 3042 25050
rect 3042 24998 3072 25050
rect 3096 24998 3106 25050
rect 3106 24998 3152 25050
rect 2856 24996 2912 24998
rect 2936 24996 2992 24998
rect 3016 24996 3072 24998
rect 3096 24996 3152 24998
rect 1356 24506 1412 24508
rect 1436 24506 1492 24508
rect 1516 24506 1572 24508
rect 1596 24506 1652 24508
rect 1356 24454 1402 24506
rect 1402 24454 1412 24506
rect 1436 24454 1466 24506
rect 1466 24454 1478 24506
rect 1478 24454 1492 24506
rect 1516 24454 1530 24506
rect 1530 24454 1542 24506
rect 1542 24454 1572 24506
rect 1596 24454 1606 24506
rect 1606 24454 1652 24506
rect 1356 24452 1412 24454
rect 1436 24452 1492 24454
rect 1516 24452 1572 24454
rect 1596 24452 1652 24454
rect 4356 24506 4412 24508
rect 4436 24506 4492 24508
rect 4516 24506 4572 24508
rect 4596 24506 4652 24508
rect 4356 24454 4402 24506
rect 4402 24454 4412 24506
rect 4436 24454 4466 24506
rect 4466 24454 4478 24506
rect 4478 24454 4492 24506
rect 4516 24454 4530 24506
rect 4530 24454 4542 24506
rect 4542 24454 4572 24506
rect 4596 24454 4606 24506
rect 4606 24454 4652 24506
rect 4356 24452 4412 24454
rect 4436 24452 4492 24454
rect 4516 24452 4572 24454
rect 4596 24452 4652 24454
rect 2856 23962 2912 23964
rect 2936 23962 2992 23964
rect 3016 23962 3072 23964
rect 3096 23962 3152 23964
rect 2856 23910 2902 23962
rect 2902 23910 2912 23962
rect 2936 23910 2966 23962
rect 2966 23910 2978 23962
rect 2978 23910 2992 23962
rect 3016 23910 3030 23962
rect 3030 23910 3042 23962
rect 3042 23910 3072 23962
rect 3096 23910 3106 23962
rect 3106 23910 3152 23962
rect 2856 23908 2912 23910
rect 2936 23908 2992 23910
rect 3016 23908 3072 23910
rect 3096 23908 3152 23910
rect 1356 23418 1412 23420
rect 1436 23418 1492 23420
rect 1516 23418 1572 23420
rect 1596 23418 1652 23420
rect 1356 23366 1402 23418
rect 1402 23366 1412 23418
rect 1436 23366 1466 23418
rect 1466 23366 1478 23418
rect 1478 23366 1492 23418
rect 1516 23366 1530 23418
rect 1530 23366 1542 23418
rect 1542 23366 1572 23418
rect 1596 23366 1606 23418
rect 1606 23366 1652 23418
rect 1356 23364 1412 23366
rect 1436 23364 1492 23366
rect 1516 23364 1572 23366
rect 1596 23364 1652 23366
rect 2856 22874 2912 22876
rect 2936 22874 2992 22876
rect 3016 22874 3072 22876
rect 3096 22874 3152 22876
rect 2856 22822 2902 22874
rect 2902 22822 2912 22874
rect 2936 22822 2966 22874
rect 2966 22822 2978 22874
rect 2978 22822 2992 22874
rect 3016 22822 3030 22874
rect 3030 22822 3042 22874
rect 3042 22822 3072 22874
rect 3096 22822 3106 22874
rect 3106 22822 3152 22874
rect 2856 22820 2912 22822
rect 2936 22820 2992 22822
rect 3016 22820 3072 22822
rect 3096 22820 3152 22822
rect 4356 23418 4412 23420
rect 4436 23418 4492 23420
rect 4516 23418 4572 23420
rect 4596 23418 4652 23420
rect 4356 23366 4402 23418
rect 4402 23366 4412 23418
rect 4436 23366 4466 23418
rect 4466 23366 4478 23418
rect 4478 23366 4492 23418
rect 4516 23366 4530 23418
rect 4530 23366 4542 23418
rect 4542 23366 4572 23418
rect 4596 23366 4606 23418
rect 4606 23366 4652 23418
rect 4356 23364 4412 23366
rect 4436 23364 4492 23366
rect 4516 23364 4572 23366
rect 4596 23364 4652 23366
rect 1356 22330 1412 22332
rect 1436 22330 1492 22332
rect 1516 22330 1572 22332
rect 1596 22330 1652 22332
rect 1356 22278 1402 22330
rect 1402 22278 1412 22330
rect 1436 22278 1466 22330
rect 1466 22278 1478 22330
rect 1478 22278 1492 22330
rect 1516 22278 1530 22330
rect 1530 22278 1542 22330
rect 1542 22278 1572 22330
rect 1596 22278 1606 22330
rect 1606 22278 1652 22330
rect 1356 22276 1412 22278
rect 1436 22276 1492 22278
rect 1516 22276 1572 22278
rect 1596 22276 1652 22278
rect 4356 22330 4412 22332
rect 4436 22330 4492 22332
rect 4516 22330 4572 22332
rect 4596 22330 4652 22332
rect 4356 22278 4402 22330
rect 4402 22278 4412 22330
rect 4436 22278 4466 22330
rect 4466 22278 4478 22330
rect 4478 22278 4492 22330
rect 4516 22278 4530 22330
rect 4530 22278 4542 22330
rect 4542 22278 4572 22330
rect 4596 22278 4606 22330
rect 4606 22278 4652 22330
rect 4356 22276 4412 22278
rect 4436 22276 4492 22278
rect 4516 22276 4572 22278
rect 4596 22276 4652 22278
rect 2856 21786 2912 21788
rect 2936 21786 2992 21788
rect 3016 21786 3072 21788
rect 3096 21786 3152 21788
rect 2856 21734 2902 21786
rect 2902 21734 2912 21786
rect 2936 21734 2966 21786
rect 2966 21734 2978 21786
rect 2978 21734 2992 21786
rect 3016 21734 3030 21786
rect 3030 21734 3042 21786
rect 3042 21734 3072 21786
rect 3096 21734 3106 21786
rect 3106 21734 3152 21786
rect 2856 21732 2912 21734
rect 2936 21732 2992 21734
rect 3016 21732 3072 21734
rect 3096 21732 3152 21734
rect 1356 21242 1412 21244
rect 1436 21242 1492 21244
rect 1516 21242 1572 21244
rect 1596 21242 1652 21244
rect 1356 21190 1402 21242
rect 1402 21190 1412 21242
rect 1436 21190 1466 21242
rect 1466 21190 1478 21242
rect 1478 21190 1492 21242
rect 1516 21190 1530 21242
rect 1530 21190 1542 21242
rect 1542 21190 1572 21242
rect 1596 21190 1606 21242
rect 1606 21190 1652 21242
rect 1356 21188 1412 21190
rect 1436 21188 1492 21190
rect 1516 21188 1572 21190
rect 1596 21188 1652 21190
rect 2856 20698 2912 20700
rect 2936 20698 2992 20700
rect 3016 20698 3072 20700
rect 3096 20698 3152 20700
rect 2856 20646 2902 20698
rect 2902 20646 2912 20698
rect 2936 20646 2966 20698
rect 2966 20646 2978 20698
rect 2978 20646 2992 20698
rect 3016 20646 3030 20698
rect 3030 20646 3042 20698
rect 3042 20646 3072 20698
rect 3096 20646 3106 20698
rect 3106 20646 3152 20698
rect 2856 20644 2912 20646
rect 2936 20644 2992 20646
rect 3016 20644 3072 20646
rect 3096 20644 3152 20646
rect 4356 21242 4412 21244
rect 4436 21242 4492 21244
rect 4516 21242 4572 21244
rect 4596 21242 4652 21244
rect 4356 21190 4402 21242
rect 4402 21190 4412 21242
rect 4436 21190 4466 21242
rect 4466 21190 4478 21242
rect 4478 21190 4492 21242
rect 4516 21190 4530 21242
rect 4530 21190 4542 21242
rect 4542 21190 4572 21242
rect 4596 21190 4606 21242
rect 4606 21190 4652 21242
rect 4356 21188 4412 21190
rect 4436 21188 4492 21190
rect 4516 21188 4572 21190
rect 4596 21188 4652 21190
rect 5856 25050 5912 25052
rect 5936 25050 5992 25052
rect 6016 25050 6072 25052
rect 6096 25050 6152 25052
rect 5856 24998 5902 25050
rect 5902 24998 5912 25050
rect 5936 24998 5966 25050
rect 5966 24998 5978 25050
rect 5978 24998 5992 25050
rect 6016 24998 6030 25050
rect 6030 24998 6042 25050
rect 6042 24998 6072 25050
rect 6096 24998 6106 25050
rect 6106 24998 6152 25050
rect 5856 24996 5912 24998
rect 5936 24996 5992 24998
rect 6016 24996 6072 24998
rect 6096 24996 6152 24998
rect 5856 23962 5912 23964
rect 5936 23962 5992 23964
rect 6016 23962 6072 23964
rect 6096 23962 6152 23964
rect 5856 23910 5902 23962
rect 5902 23910 5912 23962
rect 5936 23910 5966 23962
rect 5966 23910 5978 23962
rect 5978 23910 5992 23962
rect 6016 23910 6030 23962
rect 6030 23910 6042 23962
rect 6042 23910 6072 23962
rect 6096 23910 6106 23962
rect 6106 23910 6152 23962
rect 5856 23908 5912 23910
rect 5936 23908 5992 23910
rect 6016 23908 6072 23910
rect 6096 23908 6152 23910
rect 5170 21936 5226 21992
rect 5856 22874 5912 22876
rect 5936 22874 5992 22876
rect 6016 22874 6072 22876
rect 6096 22874 6152 22876
rect 5856 22822 5902 22874
rect 5902 22822 5912 22874
rect 5936 22822 5966 22874
rect 5966 22822 5978 22874
rect 5978 22822 5992 22874
rect 6016 22822 6030 22874
rect 6030 22822 6042 22874
rect 6042 22822 6072 22874
rect 6096 22822 6106 22874
rect 6106 22822 6152 22874
rect 5856 22820 5912 22822
rect 5936 22820 5992 22822
rect 6016 22820 6072 22822
rect 6096 22820 6152 22822
rect 1356 20154 1412 20156
rect 1436 20154 1492 20156
rect 1516 20154 1572 20156
rect 1596 20154 1652 20156
rect 1356 20102 1402 20154
rect 1402 20102 1412 20154
rect 1436 20102 1466 20154
rect 1466 20102 1478 20154
rect 1478 20102 1492 20154
rect 1516 20102 1530 20154
rect 1530 20102 1542 20154
rect 1542 20102 1572 20154
rect 1596 20102 1606 20154
rect 1606 20102 1652 20154
rect 1356 20100 1412 20102
rect 1436 20100 1492 20102
rect 1516 20100 1572 20102
rect 1596 20100 1652 20102
rect 2856 19610 2912 19612
rect 2936 19610 2992 19612
rect 3016 19610 3072 19612
rect 3096 19610 3152 19612
rect 2856 19558 2902 19610
rect 2902 19558 2912 19610
rect 2936 19558 2966 19610
rect 2966 19558 2978 19610
rect 2978 19558 2992 19610
rect 3016 19558 3030 19610
rect 3030 19558 3042 19610
rect 3042 19558 3072 19610
rect 3096 19558 3106 19610
rect 3106 19558 3152 19610
rect 2856 19556 2912 19558
rect 2936 19556 2992 19558
rect 3016 19556 3072 19558
rect 3096 19556 3152 19558
rect 1214 19116 1216 19136
rect 1216 19116 1268 19136
rect 1268 19116 1270 19136
rect 1214 19080 1270 19116
rect 1356 19066 1412 19068
rect 1436 19066 1492 19068
rect 1516 19066 1572 19068
rect 1596 19066 1652 19068
rect 1356 19014 1402 19066
rect 1402 19014 1412 19066
rect 1436 19014 1466 19066
rect 1466 19014 1478 19066
rect 1478 19014 1492 19066
rect 1516 19014 1530 19066
rect 1530 19014 1542 19066
rect 1542 19014 1572 19066
rect 1596 19014 1606 19066
rect 1606 19014 1652 19066
rect 1356 19012 1412 19014
rect 1436 19012 1492 19014
rect 1516 19012 1572 19014
rect 1596 19012 1652 19014
rect 4356 20154 4412 20156
rect 4436 20154 4492 20156
rect 4516 20154 4572 20156
rect 4596 20154 4652 20156
rect 4356 20102 4402 20154
rect 4402 20102 4412 20154
rect 4436 20102 4466 20154
rect 4466 20102 4478 20154
rect 4478 20102 4492 20154
rect 4516 20102 4530 20154
rect 4530 20102 4542 20154
rect 4542 20102 4572 20154
rect 4596 20102 4606 20154
rect 4606 20102 4652 20154
rect 4356 20100 4412 20102
rect 4436 20100 4492 20102
rect 4516 20100 4572 20102
rect 4596 20100 4652 20102
rect 5856 21786 5912 21788
rect 5936 21786 5992 21788
rect 6016 21786 6072 21788
rect 6096 21786 6152 21788
rect 5856 21734 5902 21786
rect 5902 21734 5912 21786
rect 5936 21734 5966 21786
rect 5966 21734 5978 21786
rect 5978 21734 5992 21786
rect 6016 21734 6030 21786
rect 6030 21734 6042 21786
rect 6042 21734 6072 21786
rect 6096 21734 6106 21786
rect 6106 21734 6152 21786
rect 5856 21732 5912 21734
rect 5936 21732 5992 21734
rect 6016 21732 6072 21734
rect 6096 21732 6152 21734
rect 2856 18522 2912 18524
rect 2936 18522 2992 18524
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 2856 18470 2902 18522
rect 2902 18470 2912 18522
rect 2936 18470 2966 18522
rect 2966 18470 2978 18522
rect 2978 18470 2992 18522
rect 3016 18470 3030 18522
rect 3030 18470 3042 18522
rect 3042 18470 3072 18522
rect 3096 18470 3106 18522
rect 3106 18470 3152 18522
rect 2856 18468 2912 18470
rect 2936 18468 2992 18470
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 386 18400 442 18456
rect 4356 19066 4412 19068
rect 4436 19066 4492 19068
rect 4516 19066 4572 19068
rect 4596 19066 4652 19068
rect 4356 19014 4402 19066
rect 4402 19014 4412 19066
rect 4436 19014 4466 19066
rect 4466 19014 4478 19066
rect 4478 19014 4492 19066
rect 4516 19014 4530 19066
rect 4530 19014 4542 19066
rect 4542 19014 4572 19066
rect 4596 19014 4606 19066
rect 4606 19014 4652 19066
rect 4356 19012 4412 19014
rect 4436 19012 4492 19014
rect 4516 19012 4572 19014
rect 4596 19012 4652 19014
rect 5856 20698 5912 20700
rect 5936 20698 5992 20700
rect 6016 20698 6072 20700
rect 6096 20698 6152 20700
rect 5856 20646 5902 20698
rect 5902 20646 5912 20698
rect 5936 20646 5966 20698
rect 5966 20646 5978 20698
rect 5978 20646 5992 20698
rect 6016 20646 6030 20698
rect 6030 20646 6042 20698
rect 6042 20646 6072 20698
rect 6096 20646 6106 20698
rect 6106 20646 6152 20698
rect 5856 20644 5912 20646
rect 5936 20644 5992 20646
rect 6016 20644 6072 20646
rect 6096 20644 6152 20646
rect 5856 19610 5912 19612
rect 5936 19610 5992 19612
rect 6016 19610 6072 19612
rect 6096 19610 6152 19612
rect 5856 19558 5902 19610
rect 5902 19558 5912 19610
rect 5936 19558 5966 19610
rect 5966 19558 5978 19610
rect 5978 19558 5992 19610
rect 6016 19558 6030 19610
rect 6030 19558 6042 19610
rect 6042 19558 6072 19610
rect 6096 19558 6106 19610
rect 6106 19558 6152 19610
rect 5856 19556 5912 19558
rect 5936 19556 5992 19558
rect 6016 19556 6072 19558
rect 6096 19556 6152 19558
rect 1356 17978 1412 17980
rect 1436 17978 1492 17980
rect 1516 17978 1572 17980
rect 1596 17978 1652 17980
rect 1356 17926 1402 17978
rect 1402 17926 1412 17978
rect 1436 17926 1466 17978
rect 1466 17926 1478 17978
rect 1478 17926 1492 17978
rect 1516 17926 1530 17978
rect 1530 17926 1542 17978
rect 1542 17926 1572 17978
rect 1596 17926 1606 17978
rect 1606 17926 1652 17978
rect 1356 17924 1412 17926
rect 1436 17924 1492 17926
rect 1516 17924 1572 17926
rect 1596 17924 1652 17926
rect 4356 17978 4412 17980
rect 4436 17978 4492 17980
rect 4516 17978 4572 17980
rect 4596 17978 4652 17980
rect 4356 17926 4402 17978
rect 4402 17926 4412 17978
rect 4436 17926 4466 17978
rect 4466 17926 4478 17978
rect 4478 17926 4492 17978
rect 4516 17926 4530 17978
rect 4530 17926 4542 17978
rect 4542 17926 4572 17978
rect 4596 17926 4606 17978
rect 4606 17926 4652 17978
rect 4356 17924 4412 17926
rect 4436 17924 4492 17926
rect 4516 17924 4572 17926
rect 4596 17924 4652 17926
rect 2856 17434 2912 17436
rect 2936 17434 2992 17436
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 2856 17382 2902 17434
rect 2902 17382 2912 17434
rect 2936 17382 2966 17434
rect 2966 17382 2978 17434
rect 2978 17382 2992 17434
rect 3016 17382 3030 17434
rect 3030 17382 3042 17434
rect 3042 17382 3072 17434
rect 3096 17382 3106 17434
rect 3106 17382 3152 17434
rect 2856 17380 2912 17382
rect 2936 17380 2992 17382
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 7356 24506 7412 24508
rect 7436 24506 7492 24508
rect 7516 24506 7572 24508
rect 7596 24506 7652 24508
rect 7356 24454 7402 24506
rect 7402 24454 7412 24506
rect 7436 24454 7466 24506
rect 7466 24454 7478 24506
rect 7478 24454 7492 24506
rect 7516 24454 7530 24506
rect 7530 24454 7542 24506
rect 7542 24454 7572 24506
rect 7596 24454 7606 24506
rect 7606 24454 7652 24506
rect 7356 24452 7412 24454
rect 7436 24452 7492 24454
rect 7516 24452 7572 24454
rect 7596 24452 7652 24454
rect 7356 23418 7412 23420
rect 7436 23418 7492 23420
rect 7516 23418 7572 23420
rect 7596 23418 7652 23420
rect 7356 23366 7402 23418
rect 7402 23366 7412 23418
rect 7436 23366 7466 23418
rect 7466 23366 7478 23418
rect 7478 23366 7492 23418
rect 7516 23366 7530 23418
rect 7530 23366 7542 23418
rect 7542 23366 7572 23418
rect 7596 23366 7606 23418
rect 7606 23366 7652 23418
rect 7356 23364 7412 23366
rect 7436 23364 7492 23366
rect 7516 23364 7572 23366
rect 7596 23364 7652 23366
rect 7356 22330 7412 22332
rect 7436 22330 7492 22332
rect 7516 22330 7572 22332
rect 7596 22330 7652 22332
rect 7356 22278 7402 22330
rect 7402 22278 7412 22330
rect 7436 22278 7466 22330
rect 7466 22278 7478 22330
rect 7478 22278 7492 22330
rect 7516 22278 7530 22330
rect 7530 22278 7542 22330
rect 7542 22278 7572 22330
rect 7596 22278 7606 22330
rect 7606 22278 7652 22330
rect 7356 22276 7412 22278
rect 7436 22276 7492 22278
rect 7516 22276 7572 22278
rect 7596 22276 7652 22278
rect 7654 21956 7710 21992
rect 7654 21936 7656 21956
rect 7656 21936 7708 21956
rect 7708 21936 7710 21956
rect 7356 21242 7412 21244
rect 7436 21242 7492 21244
rect 7516 21242 7572 21244
rect 7596 21242 7652 21244
rect 7356 21190 7402 21242
rect 7402 21190 7412 21242
rect 7436 21190 7466 21242
rect 7466 21190 7478 21242
rect 7478 21190 7492 21242
rect 7516 21190 7530 21242
rect 7530 21190 7542 21242
rect 7542 21190 7572 21242
rect 7596 21190 7606 21242
rect 7606 21190 7652 21242
rect 7356 21188 7412 21190
rect 7436 21188 7492 21190
rect 7516 21188 7572 21190
rect 7596 21188 7652 21190
rect 7356 20154 7412 20156
rect 7436 20154 7492 20156
rect 7516 20154 7572 20156
rect 7596 20154 7652 20156
rect 7356 20102 7402 20154
rect 7402 20102 7412 20154
rect 7436 20102 7466 20154
rect 7466 20102 7478 20154
rect 7478 20102 7492 20154
rect 7516 20102 7530 20154
rect 7530 20102 7542 20154
rect 7542 20102 7572 20154
rect 7596 20102 7606 20154
rect 7606 20102 7652 20154
rect 7356 20100 7412 20102
rect 7436 20100 7492 20102
rect 7516 20100 7572 20102
rect 7596 20100 7652 20102
rect 5856 18522 5912 18524
rect 5936 18522 5992 18524
rect 6016 18522 6072 18524
rect 6096 18522 6152 18524
rect 5856 18470 5902 18522
rect 5902 18470 5912 18522
rect 5936 18470 5966 18522
rect 5966 18470 5978 18522
rect 5978 18470 5992 18522
rect 6016 18470 6030 18522
rect 6030 18470 6042 18522
rect 6042 18470 6072 18522
rect 6096 18470 6106 18522
rect 6106 18470 6152 18522
rect 5856 18468 5912 18470
rect 5936 18468 5992 18470
rect 6016 18468 6072 18470
rect 6096 18468 6152 18470
rect 5856 17434 5912 17436
rect 5936 17434 5992 17436
rect 6016 17434 6072 17436
rect 6096 17434 6152 17436
rect 5856 17382 5902 17434
rect 5902 17382 5912 17434
rect 5936 17382 5966 17434
rect 5966 17382 5978 17434
rect 5978 17382 5992 17434
rect 6016 17382 6030 17434
rect 6030 17382 6042 17434
rect 6042 17382 6072 17434
rect 6096 17382 6106 17434
rect 6106 17382 6152 17434
rect 5856 17380 5912 17382
rect 5936 17380 5992 17382
rect 6016 17380 6072 17382
rect 6096 17380 6152 17382
rect 1356 16890 1412 16892
rect 1436 16890 1492 16892
rect 1516 16890 1572 16892
rect 1596 16890 1652 16892
rect 1356 16838 1402 16890
rect 1402 16838 1412 16890
rect 1436 16838 1466 16890
rect 1466 16838 1478 16890
rect 1478 16838 1492 16890
rect 1516 16838 1530 16890
rect 1530 16838 1542 16890
rect 1542 16838 1572 16890
rect 1596 16838 1606 16890
rect 1606 16838 1652 16890
rect 1356 16836 1412 16838
rect 1436 16836 1492 16838
rect 1516 16836 1572 16838
rect 1596 16836 1652 16838
rect 1306 16396 1308 16416
rect 1308 16396 1360 16416
rect 1360 16396 1362 16416
rect 1306 16360 1362 16396
rect 2856 16346 2912 16348
rect 2936 16346 2992 16348
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 2856 16294 2902 16346
rect 2902 16294 2912 16346
rect 2936 16294 2966 16346
rect 2966 16294 2978 16346
rect 2978 16294 2992 16346
rect 3016 16294 3030 16346
rect 3030 16294 3042 16346
rect 3042 16294 3072 16346
rect 3096 16294 3106 16346
rect 3106 16294 3152 16346
rect 2856 16292 2912 16294
rect 2936 16292 2992 16294
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 4356 16890 4412 16892
rect 4436 16890 4492 16892
rect 4516 16890 4572 16892
rect 4596 16890 4652 16892
rect 4356 16838 4402 16890
rect 4402 16838 4412 16890
rect 4436 16838 4466 16890
rect 4466 16838 4478 16890
rect 4478 16838 4492 16890
rect 4516 16838 4530 16890
rect 4530 16838 4542 16890
rect 4542 16838 4572 16890
rect 4596 16838 4606 16890
rect 4606 16838 4652 16890
rect 4356 16836 4412 16838
rect 4436 16836 4492 16838
rect 4516 16836 4572 16838
rect 4596 16836 4652 16838
rect 1356 15802 1412 15804
rect 1436 15802 1492 15804
rect 1516 15802 1572 15804
rect 1596 15802 1652 15804
rect 1356 15750 1402 15802
rect 1402 15750 1412 15802
rect 1436 15750 1466 15802
rect 1466 15750 1478 15802
rect 1478 15750 1492 15802
rect 1516 15750 1530 15802
rect 1530 15750 1542 15802
rect 1542 15750 1572 15802
rect 1596 15750 1606 15802
rect 1606 15750 1652 15802
rect 1356 15748 1412 15750
rect 1436 15748 1492 15750
rect 1516 15748 1572 15750
rect 1596 15748 1652 15750
rect 754 15680 810 15736
rect 1398 15000 1454 15056
rect 754 14320 810 14376
rect 1356 14714 1412 14716
rect 1436 14714 1492 14716
rect 1516 14714 1572 14716
rect 1596 14714 1652 14716
rect 1356 14662 1402 14714
rect 1402 14662 1412 14714
rect 1436 14662 1466 14714
rect 1466 14662 1478 14714
rect 1478 14662 1492 14714
rect 1516 14662 1530 14714
rect 1530 14662 1542 14714
rect 1542 14662 1572 14714
rect 1596 14662 1606 14714
rect 1606 14662 1652 14714
rect 1356 14660 1412 14662
rect 1436 14660 1492 14662
rect 1516 14660 1572 14662
rect 1596 14660 1652 14662
rect 1214 13640 1270 13696
rect 1356 13626 1412 13628
rect 1436 13626 1492 13628
rect 1516 13626 1572 13628
rect 1596 13626 1652 13628
rect 1356 13574 1402 13626
rect 1402 13574 1412 13626
rect 1436 13574 1466 13626
rect 1466 13574 1478 13626
rect 1478 13574 1492 13626
rect 1516 13574 1530 13626
rect 1530 13574 1542 13626
rect 1542 13574 1572 13626
rect 1596 13574 1606 13626
rect 1606 13574 1652 13626
rect 1356 13572 1412 13574
rect 1436 13572 1492 13574
rect 1516 13572 1572 13574
rect 1596 13572 1652 13574
rect 1306 12980 1362 13016
rect 1306 12960 1308 12980
rect 1308 12960 1360 12980
rect 1360 12960 1362 12980
rect 2856 15258 2912 15260
rect 2936 15258 2992 15260
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 2856 15206 2902 15258
rect 2902 15206 2912 15258
rect 2936 15206 2966 15258
rect 2966 15206 2978 15258
rect 2978 15206 2992 15258
rect 3016 15206 3030 15258
rect 3030 15206 3042 15258
rect 3042 15206 3072 15258
rect 3096 15206 3106 15258
rect 3106 15206 3152 15258
rect 2856 15204 2912 15206
rect 2936 15204 2992 15206
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 4356 15802 4412 15804
rect 4436 15802 4492 15804
rect 4516 15802 4572 15804
rect 4596 15802 4652 15804
rect 4356 15750 4402 15802
rect 4402 15750 4412 15802
rect 4436 15750 4466 15802
rect 4466 15750 4478 15802
rect 4478 15750 4492 15802
rect 4516 15750 4530 15802
rect 4530 15750 4542 15802
rect 4542 15750 4572 15802
rect 4596 15750 4606 15802
rect 4606 15750 4652 15802
rect 4356 15748 4412 15750
rect 4436 15748 4492 15750
rect 4516 15748 4572 15750
rect 4596 15748 4652 15750
rect 7356 19066 7412 19068
rect 7436 19066 7492 19068
rect 7516 19066 7572 19068
rect 7596 19066 7652 19068
rect 7356 19014 7402 19066
rect 7402 19014 7412 19066
rect 7436 19014 7466 19066
rect 7466 19014 7478 19066
rect 7478 19014 7492 19066
rect 7516 19014 7530 19066
rect 7530 19014 7542 19066
rect 7542 19014 7572 19066
rect 7596 19014 7606 19066
rect 7606 19014 7652 19066
rect 7356 19012 7412 19014
rect 7436 19012 7492 19014
rect 7516 19012 7572 19014
rect 7596 19012 7652 19014
rect 8856 25050 8912 25052
rect 8936 25050 8992 25052
rect 9016 25050 9072 25052
rect 9096 25050 9152 25052
rect 8856 24998 8902 25050
rect 8902 24998 8912 25050
rect 8936 24998 8966 25050
rect 8966 24998 8978 25050
rect 8978 24998 8992 25050
rect 9016 24998 9030 25050
rect 9030 24998 9042 25050
rect 9042 24998 9072 25050
rect 9096 24998 9106 25050
rect 9106 24998 9152 25050
rect 8856 24996 8912 24998
rect 8936 24996 8992 24998
rect 9016 24996 9072 24998
rect 9096 24996 9152 24998
rect 8856 23962 8912 23964
rect 8936 23962 8992 23964
rect 9016 23962 9072 23964
rect 9096 23962 9152 23964
rect 8856 23910 8902 23962
rect 8902 23910 8912 23962
rect 8936 23910 8966 23962
rect 8966 23910 8978 23962
rect 8978 23910 8992 23962
rect 9016 23910 9030 23962
rect 9030 23910 9042 23962
rect 9042 23910 9072 23962
rect 9096 23910 9106 23962
rect 9106 23910 9152 23962
rect 8856 23908 8912 23910
rect 8936 23908 8992 23910
rect 9016 23908 9072 23910
rect 9096 23908 9152 23910
rect 8856 22874 8912 22876
rect 8936 22874 8992 22876
rect 9016 22874 9072 22876
rect 9096 22874 9152 22876
rect 8856 22822 8902 22874
rect 8902 22822 8912 22874
rect 8936 22822 8966 22874
rect 8966 22822 8978 22874
rect 8978 22822 8992 22874
rect 9016 22822 9030 22874
rect 9030 22822 9042 22874
rect 9042 22822 9072 22874
rect 9096 22822 9106 22874
rect 9106 22822 9152 22874
rect 8856 22820 8912 22822
rect 8936 22820 8992 22822
rect 9016 22820 9072 22822
rect 9096 22820 9152 22822
rect 10356 24506 10412 24508
rect 10436 24506 10492 24508
rect 10516 24506 10572 24508
rect 10596 24506 10652 24508
rect 10356 24454 10402 24506
rect 10402 24454 10412 24506
rect 10436 24454 10466 24506
rect 10466 24454 10478 24506
rect 10478 24454 10492 24506
rect 10516 24454 10530 24506
rect 10530 24454 10542 24506
rect 10542 24454 10572 24506
rect 10596 24454 10606 24506
rect 10606 24454 10652 24506
rect 10356 24452 10412 24454
rect 10436 24452 10492 24454
rect 10516 24452 10572 24454
rect 10596 24452 10652 24454
rect 10356 23418 10412 23420
rect 10436 23418 10492 23420
rect 10516 23418 10572 23420
rect 10596 23418 10652 23420
rect 10356 23366 10402 23418
rect 10402 23366 10412 23418
rect 10436 23366 10466 23418
rect 10466 23366 10478 23418
rect 10478 23366 10492 23418
rect 10516 23366 10530 23418
rect 10530 23366 10542 23418
rect 10542 23366 10572 23418
rect 10596 23366 10606 23418
rect 10606 23366 10652 23418
rect 10356 23364 10412 23366
rect 10436 23364 10492 23366
rect 10516 23364 10572 23366
rect 10596 23364 10652 23366
rect 8856 21786 8912 21788
rect 8936 21786 8992 21788
rect 9016 21786 9072 21788
rect 9096 21786 9152 21788
rect 8856 21734 8902 21786
rect 8902 21734 8912 21786
rect 8936 21734 8966 21786
rect 8966 21734 8978 21786
rect 8978 21734 8992 21786
rect 9016 21734 9030 21786
rect 9030 21734 9042 21786
rect 9042 21734 9072 21786
rect 9096 21734 9106 21786
rect 9106 21734 9152 21786
rect 8856 21732 8912 21734
rect 8936 21732 8992 21734
rect 9016 21732 9072 21734
rect 9096 21732 9152 21734
rect 8856 20698 8912 20700
rect 8936 20698 8992 20700
rect 9016 20698 9072 20700
rect 9096 20698 9152 20700
rect 8856 20646 8902 20698
rect 8902 20646 8912 20698
rect 8936 20646 8966 20698
rect 8966 20646 8978 20698
rect 8978 20646 8992 20698
rect 9016 20646 9030 20698
rect 9030 20646 9042 20698
rect 9042 20646 9072 20698
rect 9096 20646 9106 20698
rect 9106 20646 9152 20698
rect 8856 20644 8912 20646
rect 8936 20644 8992 20646
rect 9016 20644 9072 20646
rect 9096 20644 9152 20646
rect 8856 19610 8912 19612
rect 8936 19610 8992 19612
rect 9016 19610 9072 19612
rect 9096 19610 9152 19612
rect 8856 19558 8902 19610
rect 8902 19558 8912 19610
rect 8936 19558 8966 19610
rect 8966 19558 8978 19610
rect 8978 19558 8992 19610
rect 9016 19558 9030 19610
rect 9030 19558 9042 19610
rect 9042 19558 9072 19610
rect 9096 19558 9106 19610
rect 9106 19558 9152 19610
rect 8856 19556 8912 19558
rect 8936 19556 8992 19558
rect 9016 19556 9072 19558
rect 9096 19556 9152 19558
rect 10356 22330 10412 22332
rect 10436 22330 10492 22332
rect 10516 22330 10572 22332
rect 10596 22330 10652 22332
rect 10356 22278 10402 22330
rect 10402 22278 10412 22330
rect 10436 22278 10466 22330
rect 10466 22278 10478 22330
rect 10478 22278 10492 22330
rect 10516 22278 10530 22330
rect 10530 22278 10542 22330
rect 10542 22278 10572 22330
rect 10596 22278 10606 22330
rect 10606 22278 10652 22330
rect 10356 22276 10412 22278
rect 10436 22276 10492 22278
rect 10516 22276 10572 22278
rect 10596 22276 10652 22278
rect 10356 21242 10412 21244
rect 10436 21242 10492 21244
rect 10516 21242 10572 21244
rect 10596 21242 10652 21244
rect 10356 21190 10402 21242
rect 10402 21190 10412 21242
rect 10436 21190 10466 21242
rect 10466 21190 10478 21242
rect 10478 21190 10492 21242
rect 10516 21190 10530 21242
rect 10530 21190 10542 21242
rect 10542 21190 10572 21242
rect 10596 21190 10606 21242
rect 10606 21190 10652 21242
rect 10356 21188 10412 21190
rect 10436 21188 10492 21190
rect 10516 21188 10572 21190
rect 10596 21188 10652 21190
rect 7356 17978 7412 17980
rect 7436 17978 7492 17980
rect 7516 17978 7572 17980
rect 7596 17978 7652 17980
rect 7356 17926 7402 17978
rect 7402 17926 7412 17978
rect 7436 17926 7466 17978
rect 7466 17926 7478 17978
rect 7478 17926 7492 17978
rect 7516 17926 7530 17978
rect 7530 17926 7542 17978
rect 7542 17926 7572 17978
rect 7596 17926 7606 17978
rect 7606 17926 7652 17978
rect 7356 17924 7412 17926
rect 7436 17924 7492 17926
rect 7516 17924 7572 17926
rect 7596 17924 7652 17926
rect 8856 18522 8912 18524
rect 8936 18522 8992 18524
rect 9016 18522 9072 18524
rect 9096 18522 9152 18524
rect 8856 18470 8902 18522
rect 8902 18470 8912 18522
rect 8936 18470 8966 18522
rect 8966 18470 8978 18522
rect 8978 18470 8992 18522
rect 9016 18470 9030 18522
rect 9030 18470 9042 18522
rect 9042 18470 9072 18522
rect 9096 18470 9106 18522
rect 9106 18470 9152 18522
rect 8856 18468 8912 18470
rect 8936 18468 8992 18470
rect 9016 18468 9072 18470
rect 9096 18468 9152 18470
rect 7356 16890 7412 16892
rect 7436 16890 7492 16892
rect 7516 16890 7572 16892
rect 7596 16890 7652 16892
rect 7356 16838 7402 16890
rect 7402 16838 7412 16890
rect 7436 16838 7466 16890
rect 7466 16838 7478 16890
rect 7478 16838 7492 16890
rect 7516 16838 7530 16890
rect 7530 16838 7542 16890
rect 7542 16838 7572 16890
rect 7596 16838 7606 16890
rect 7606 16838 7652 16890
rect 7356 16836 7412 16838
rect 7436 16836 7492 16838
rect 7516 16836 7572 16838
rect 7596 16836 7652 16838
rect 5856 16346 5912 16348
rect 5936 16346 5992 16348
rect 6016 16346 6072 16348
rect 6096 16346 6152 16348
rect 5856 16294 5902 16346
rect 5902 16294 5912 16346
rect 5936 16294 5966 16346
rect 5966 16294 5978 16346
rect 5978 16294 5992 16346
rect 6016 16294 6030 16346
rect 6030 16294 6042 16346
rect 6042 16294 6072 16346
rect 6096 16294 6106 16346
rect 6106 16294 6152 16346
rect 5856 16292 5912 16294
rect 5936 16292 5992 16294
rect 6016 16292 6072 16294
rect 6096 16292 6152 16294
rect 8856 17434 8912 17436
rect 8936 17434 8992 17436
rect 9016 17434 9072 17436
rect 9096 17434 9152 17436
rect 8856 17382 8902 17434
rect 8902 17382 8912 17434
rect 8936 17382 8966 17434
rect 8966 17382 8978 17434
rect 8978 17382 8992 17434
rect 9016 17382 9030 17434
rect 9030 17382 9042 17434
rect 9042 17382 9072 17434
rect 9096 17382 9106 17434
rect 9106 17382 9152 17434
rect 8856 17380 8912 17382
rect 8936 17380 8992 17382
rect 9016 17380 9072 17382
rect 9096 17380 9152 17382
rect 10356 20154 10412 20156
rect 10436 20154 10492 20156
rect 10516 20154 10572 20156
rect 10596 20154 10652 20156
rect 10356 20102 10402 20154
rect 10402 20102 10412 20154
rect 10436 20102 10466 20154
rect 10466 20102 10478 20154
rect 10478 20102 10492 20154
rect 10516 20102 10530 20154
rect 10530 20102 10542 20154
rect 10542 20102 10572 20154
rect 10596 20102 10606 20154
rect 10606 20102 10652 20154
rect 10356 20100 10412 20102
rect 10436 20100 10492 20102
rect 10516 20100 10572 20102
rect 10596 20100 10652 20102
rect 11242 23568 11298 23624
rect 11856 25050 11912 25052
rect 11936 25050 11992 25052
rect 12016 25050 12072 25052
rect 12096 25050 12152 25052
rect 11856 24998 11902 25050
rect 11902 24998 11912 25050
rect 11936 24998 11966 25050
rect 11966 24998 11978 25050
rect 11978 24998 11992 25050
rect 12016 24998 12030 25050
rect 12030 24998 12042 25050
rect 12042 24998 12072 25050
rect 12096 24998 12106 25050
rect 12106 24998 12152 25050
rect 11856 24996 11912 24998
rect 11936 24996 11992 24998
rect 12016 24996 12072 24998
rect 12096 24996 12152 24998
rect 11242 21936 11298 21992
rect 10356 19066 10412 19068
rect 10436 19066 10492 19068
rect 10516 19066 10572 19068
rect 10596 19066 10652 19068
rect 10356 19014 10402 19066
rect 10402 19014 10412 19066
rect 10436 19014 10466 19066
rect 10466 19014 10478 19066
rect 10478 19014 10492 19066
rect 10516 19014 10530 19066
rect 10530 19014 10542 19066
rect 10542 19014 10572 19066
rect 10596 19014 10606 19066
rect 10606 19014 10652 19066
rect 10356 19012 10412 19014
rect 10436 19012 10492 19014
rect 10516 19012 10572 19014
rect 10596 19012 10652 19014
rect 10356 17978 10412 17980
rect 10436 17978 10492 17980
rect 10516 17978 10572 17980
rect 10596 17978 10652 17980
rect 10356 17926 10402 17978
rect 10402 17926 10412 17978
rect 10436 17926 10466 17978
rect 10466 17926 10478 17978
rect 10478 17926 10492 17978
rect 10516 17926 10530 17978
rect 10530 17926 10542 17978
rect 10542 17926 10572 17978
rect 10596 17926 10606 17978
rect 10606 17926 10652 17978
rect 10356 17924 10412 17926
rect 10436 17924 10492 17926
rect 10516 17924 10572 17926
rect 10596 17924 10652 17926
rect 10966 18264 11022 18320
rect 8856 16346 8912 16348
rect 8936 16346 8992 16348
rect 9016 16346 9072 16348
rect 9096 16346 9152 16348
rect 8856 16294 8902 16346
rect 8902 16294 8912 16346
rect 8936 16294 8966 16346
rect 8966 16294 8978 16346
rect 8978 16294 8992 16346
rect 9016 16294 9030 16346
rect 9030 16294 9042 16346
rect 9042 16294 9072 16346
rect 9096 16294 9106 16346
rect 9106 16294 9152 16346
rect 8856 16292 8912 16294
rect 8936 16292 8992 16294
rect 9016 16292 9072 16294
rect 9096 16292 9152 16294
rect 5856 15258 5912 15260
rect 5936 15258 5992 15260
rect 6016 15258 6072 15260
rect 6096 15258 6152 15260
rect 5856 15206 5902 15258
rect 5902 15206 5912 15258
rect 5936 15206 5966 15258
rect 5966 15206 5978 15258
rect 5978 15206 5992 15258
rect 6016 15206 6030 15258
rect 6030 15206 6042 15258
rect 6042 15206 6072 15258
rect 6096 15206 6106 15258
rect 6106 15206 6152 15258
rect 5856 15204 5912 15206
rect 5936 15204 5992 15206
rect 6016 15204 6072 15206
rect 6096 15204 6152 15206
rect 2856 14170 2912 14172
rect 2936 14170 2992 14172
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 2856 14118 2902 14170
rect 2902 14118 2912 14170
rect 2936 14118 2966 14170
rect 2966 14118 2978 14170
rect 2978 14118 2992 14170
rect 3016 14118 3030 14170
rect 3030 14118 3042 14170
rect 3042 14118 3072 14170
rect 3096 14118 3106 14170
rect 3106 14118 3152 14170
rect 2856 14116 2912 14118
rect 2936 14116 2992 14118
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 2856 13082 2912 13084
rect 2936 13082 2992 13084
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 2856 13030 2902 13082
rect 2902 13030 2912 13082
rect 2936 13030 2966 13082
rect 2966 13030 2978 13082
rect 2978 13030 2992 13082
rect 3016 13030 3030 13082
rect 3030 13030 3042 13082
rect 3042 13030 3072 13082
rect 3096 13030 3106 13082
rect 3106 13030 3152 13082
rect 2856 13028 2912 13030
rect 2936 13028 2992 13030
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 1356 12538 1412 12540
rect 1436 12538 1492 12540
rect 1516 12538 1572 12540
rect 1596 12538 1652 12540
rect 1356 12486 1402 12538
rect 1402 12486 1412 12538
rect 1436 12486 1466 12538
rect 1466 12486 1478 12538
rect 1478 12486 1492 12538
rect 1516 12486 1530 12538
rect 1530 12486 1542 12538
rect 1542 12486 1572 12538
rect 1596 12486 1606 12538
rect 1606 12486 1652 12538
rect 1356 12484 1412 12486
rect 1436 12484 1492 12486
rect 1516 12484 1572 12486
rect 1596 12484 1652 12486
rect 386 12280 442 12336
rect 2856 11994 2912 11996
rect 2936 11994 2992 11996
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 2856 11942 2902 11994
rect 2902 11942 2912 11994
rect 2936 11942 2966 11994
rect 2966 11942 2978 11994
rect 2978 11942 2992 11994
rect 3016 11942 3030 11994
rect 3030 11942 3042 11994
rect 3042 11942 3072 11994
rect 3096 11942 3106 11994
rect 3106 11942 3152 11994
rect 2856 11940 2912 11942
rect 2936 11940 2992 11942
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 4356 14714 4412 14716
rect 4436 14714 4492 14716
rect 4516 14714 4572 14716
rect 4596 14714 4652 14716
rect 4356 14662 4402 14714
rect 4402 14662 4412 14714
rect 4436 14662 4466 14714
rect 4466 14662 4478 14714
rect 4478 14662 4492 14714
rect 4516 14662 4530 14714
rect 4530 14662 4542 14714
rect 4542 14662 4572 14714
rect 4596 14662 4606 14714
rect 4606 14662 4652 14714
rect 4356 14660 4412 14662
rect 4436 14660 4492 14662
rect 4516 14660 4572 14662
rect 4596 14660 4652 14662
rect 7356 15802 7412 15804
rect 7436 15802 7492 15804
rect 7516 15802 7572 15804
rect 7596 15802 7652 15804
rect 7356 15750 7402 15802
rect 7402 15750 7412 15802
rect 7436 15750 7466 15802
rect 7466 15750 7478 15802
rect 7478 15750 7492 15802
rect 7516 15750 7530 15802
rect 7530 15750 7542 15802
rect 7542 15750 7572 15802
rect 7596 15750 7606 15802
rect 7606 15750 7652 15802
rect 7356 15748 7412 15750
rect 7436 15748 7492 15750
rect 7516 15748 7572 15750
rect 7596 15748 7652 15750
rect 4356 13626 4412 13628
rect 4436 13626 4492 13628
rect 4516 13626 4572 13628
rect 4596 13626 4652 13628
rect 4356 13574 4402 13626
rect 4402 13574 4412 13626
rect 4436 13574 4466 13626
rect 4466 13574 4478 13626
rect 4478 13574 4492 13626
rect 4516 13574 4530 13626
rect 4530 13574 4542 13626
rect 4542 13574 4572 13626
rect 4596 13574 4606 13626
rect 4606 13574 4652 13626
rect 4356 13572 4412 13574
rect 4436 13572 4492 13574
rect 4516 13572 4572 13574
rect 4596 13572 4652 13574
rect 3882 12688 3938 12744
rect 386 11600 442 11656
rect 1356 11450 1412 11452
rect 1436 11450 1492 11452
rect 1516 11450 1572 11452
rect 1596 11450 1652 11452
rect 1356 11398 1402 11450
rect 1402 11398 1412 11450
rect 1436 11398 1466 11450
rect 1466 11398 1478 11450
rect 1478 11398 1492 11450
rect 1516 11398 1530 11450
rect 1530 11398 1542 11450
rect 1542 11398 1572 11450
rect 1596 11398 1606 11450
rect 1606 11398 1652 11450
rect 1356 11396 1412 11398
rect 1436 11396 1492 11398
rect 1516 11396 1572 11398
rect 1596 11396 1652 11398
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 2856 10906 2912 10908
rect 2936 10906 2992 10908
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 2856 10854 2902 10906
rect 2902 10854 2912 10906
rect 2936 10854 2966 10906
rect 2966 10854 2978 10906
rect 2978 10854 2992 10906
rect 3016 10854 3030 10906
rect 3030 10854 3042 10906
rect 3042 10854 3072 10906
rect 3096 10854 3106 10906
rect 3106 10854 3152 10906
rect 2856 10852 2912 10854
rect 2936 10852 2992 10854
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 1858 10512 1914 10568
rect 1356 10362 1412 10364
rect 1436 10362 1492 10364
rect 1516 10362 1572 10364
rect 1596 10362 1652 10364
rect 1356 10310 1402 10362
rect 1402 10310 1412 10362
rect 1436 10310 1466 10362
rect 1466 10310 1478 10362
rect 1478 10310 1492 10362
rect 1516 10310 1530 10362
rect 1530 10310 1542 10362
rect 1542 10310 1572 10362
rect 1596 10310 1606 10362
rect 1606 10310 1652 10362
rect 1356 10308 1412 10310
rect 1436 10308 1492 10310
rect 1516 10308 1572 10310
rect 1596 10308 1652 10310
rect 386 9580 442 9616
rect 386 9560 388 9580
rect 388 9560 440 9580
rect 440 9560 442 9580
rect 1356 9274 1412 9276
rect 1436 9274 1492 9276
rect 1516 9274 1572 9276
rect 1596 9274 1652 9276
rect 1356 9222 1402 9274
rect 1402 9222 1412 9274
rect 1436 9222 1466 9274
rect 1466 9222 1478 9274
rect 1478 9222 1492 9274
rect 1516 9222 1530 9274
rect 1530 9222 1542 9274
rect 1542 9222 1572 9274
rect 1596 9222 1606 9274
rect 1606 9222 1652 9274
rect 1356 9220 1412 9222
rect 1436 9220 1492 9222
rect 1516 9220 1572 9222
rect 1596 9220 1652 9222
rect 386 8916 388 8936
rect 388 8916 440 8936
rect 440 8916 442 8936
rect 386 8880 442 8916
rect 2856 9818 2912 9820
rect 2936 9818 2992 9820
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 2856 9766 2902 9818
rect 2902 9766 2912 9818
rect 2936 9766 2966 9818
rect 2966 9766 2978 9818
rect 2978 9766 2992 9818
rect 3016 9766 3030 9818
rect 3030 9766 3042 9818
rect 3042 9766 3072 9818
rect 3096 9766 3106 9818
rect 3106 9766 3152 9818
rect 2856 9764 2912 9766
rect 2936 9764 2992 9766
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 1214 8200 1270 8256
rect 1356 8186 1412 8188
rect 1436 8186 1492 8188
rect 1516 8186 1572 8188
rect 1596 8186 1652 8188
rect 1356 8134 1402 8186
rect 1402 8134 1412 8186
rect 1436 8134 1466 8186
rect 1466 8134 1478 8186
rect 1478 8134 1492 8186
rect 1516 8134 1530 8186
rect 1530 8134 1542 8186
rect 1542 8134 1572 8186
rect 1596 8134 1606 8186
rect 1606 8134 1652 8186
rect 1356 8132 1412 8134
rect 1436 8132 1492 8134
rect 1516 8132 1572 8134
rect 1596 8132 1652 8134
rect 4356 12538 4412 12540
rect 4436 12538 4492 12540
rect 4516 12538 4572 12540
rect 4596 12538 4652 12540
rect 4356 12486 4402 12538
rect 4402 12486 4412 12538
rect 4436 12486 4466 12538
rect 4466 12486 4478 12538
rect 4478 12486 4492 12538
rect 4516 12486 4530 12538
rect 4530 12486 4542 12538
rect 4542 12486 4572 12538
rect 4596 12486 4606 12538
rect 4606 12486 4652 12538
rect 4356 12484 4412 12486
rect 4436 12484 4492 12486
rect 4516 12484 4572 12486
rect 4596 12484 4652 12486
rect 4356 11450 4412 11452
rect 4436 11450 4492 11452
rect 4516 11450 4572 11452
rect 4596 11450 4652 11452
rect 4356 11398 4402 11450
rect 4402 11398 4412 11450
rect 4436 11398 4466 11450
rect 4466 11398 4478 11450
rect 4478 11398 4492 11450
rect 4516 11398 4530 11450
rect 4530 11398 4542 11450
rect 4542 11398 4572 11450
rect 4596 11398 4606 11450
rect 4606 11398 4652 11450
rect 4356 11396 4412 11398
rect 4436 11396 4492 11398
rect 4516 11396 4572 11398
rect 4596 11396 4652 11398
rect 4356 10362 4412 10364
rect 4436 10362 4492 10364
rect 4516 10362 4572 10364
rect 4596 10362 4652 10364
rect 4356 10310 4402 10362
rect 4402 10310 4412 10362
rect 4436 10310 4466 10362
rect 4466 10310 4478 10362
rect 4478 10310 4492 10362
rect 4516 10310 4530 10362
rect 4530 10310 4542 10362
rect 4542 10310 4572 10362
rect 4596 10310 4606 10362
rect 4606 10310 4652 10362
rect 4356 10308 4412 10310
rect 4436 10308 4492 10310
rect 4516 10308 4572 10310
rect 4596 10308 4652 10310
rect 4356 9274 4412 9276
rect 4436 9274 4492 9276
rect 4516 9274 4572 9276
rect 4596 9274 4652 9276
rect 4356 9222 4402 9274
rect 4402 9222 4412 9274
rect 4436 9222 4466 9274
rect 4466 9222 4478 9274
rect 4478 9222 4492 9274
rect 4516 9222 4530 9274
rect 4530 9222 4542 9274
rect 4542 9222 4572 9274
rect 4596 9222 4606 9274
rect 4606 9222 4652 9274
rect 4356 9220 4412 9222
rect 4436 9220 4492 9222
rect 4516 9220 4572 9222
rect 4596 9220 4652 9222
rect 2856 8730 2912 8732
rect 2936 8730 2992 8732
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 2856 8678 2902 8730
rect 2902 8678 2912 8730
rect 2936 8678 2966 8730
rect 2966 8678 2978 8730
rect 2978 8678 2992 8730
rect 3016 8678 3030 8730
rect 3030 8678 3042 8730
rect 3042 8678 3072 8730
rect 3096 8678 3106 8730
rect 3106 8678 3152 8730
rect 2856 8676 2912 8678
rect 2936 8676 2992 8678
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 2856 7642 2912 7644
rect 2936 7642 2992 7644
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 2856 7590 2902 7642
rect 2902 7590 2912 7642
rect 2936 7590 2966 7642
rect 2966 7590 2978 7642
rect 2978 7590 2992 7642
rect 3016 7590 3030 7642
rect 3030 7590 3042 7642
rect 3042 7590 3072 7642
rect 3096 7590 3106 7642
rect 3106 7590 3152 7642
rect 2856 7588 2912 7590
rect 2936 7588 2992 7590
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 5856 14170 5912 14172
rect 5936 14170 5992 14172
rect 6016 14170 6072 14172
rect 6096 14170 6152 14172
rect 5856 14118 5902 14170
rect 5902 14118 5912 14170
rect 5936 14118 5966 14170
rect 5966 14118 5978 14170
rect 5978 14118 5992 14170
rect 6016 14118 6030 14170
rect 6030 14118 6042 14170
rect 6042 14118 6072 14170
rect 6096 14118 6106 14170
rect 6106 14118 6152 14170
rect 5856 14116 5912 14118
rect 5936 14116 5992 14118
rect 6016 14116 6072 14118
rect 6096 14116 6152 14118
rect 7356 14714 7412 14716
rect 7436 14714 7492 14716
rect 7516 14714 7572 14716
rect 7596 14714 7652 14716
rect 7356 14662 7402 14714
rect 7402 14662 7412 14714
rect 7436 14662 7466 14714
rect 7466 14662 7478 14714
rect 7478 14662 7492 14714
rect 7516 14662 7530 14714
rect 7530 14662 7542 14714
rect 7542 14662 7572 14714
rect 7596 14662 7606 14714
rect 7606 14662 7652 14714
rect 7356 14660 7412 14662
rect 7436 14660 7492 14662
rect 7516 14660 7572 14662
rect 7596 14660 7652 14662
rect 7356 13626 7412 13628
rect 7436 13626 7492 13628
rect 7516 13626 7572 13628
rect 7596 13626 7652 13628
rect 7356 13574 7402 13626
rect 7402 13574 7412 13626
rect 7436 13574 7466 13626
rect 7466 13574 7478 13626
rect 7478 13574 7492 13626
rect 7516 13574 7530 13626
rect 7530 13574 7542 13626
rect 7542 13574 7572 13626
rect 7596 13574 7606 13626
rect 7606 13574 7652 13626
rect 7356 13572 7412 13574
rect 7436 13572 7492 13574
rect 7516 13572 7572 13574
rect 7596 13572 7652 13574
rect 10356 16890 10412 16892
rect 10436 16890 10492 16892
rect 10516 16890 10572 16892
rect 10596 16890 10652 16892
rect 10356 16838 10402 16890
rect 10402 16838 10412 16890
rect 10436 16838 10466 16890
rect 10466 16838 10478 16890
rect 10478 16838 10492 16890
rect 10516 16838 10530 16890
rect 10530 16838 10542 16890
rect 10542 16838 10572 16890
rect 10596 16838 10606 16890
rect 10606 16838 10652 16890
rect 10356 16836 10412 16838
rect 10436 16836 10492 16838
rect 10516 16836 10572 16838
rect 10596 16836 10652 16838
rect 10356 15802 10412 15804
rect 10436 15802 10492 15804
rect 10516 15802 10572 15804
rect 10596 15802 10652 15804
rect 10356 15750 10402 15802
rect 10402 15750 10412 15802
rect 10436 15750 10466 15802
rect 10466 15750 10478 15802
rect 10478 15750 10492 15802
rect 10516 15750 10530 15802
rect 10530 15750 10542 15802
rect 10542 15750 10572 15802
rect 10596 15750 10606 15802
rect 10606 15750 10652 15802
rect 10356 15748 10412 15750
rect 10436 15748 10492 15750
rect 10516 15748 10572 15750
rect 10596 15748 10652 15750
rect 8856 15258 8912 15260
rect 8936 15258 8992 15260
rect 9016 15258 9072 15260
rect 9096 15258 9152 15260
rect 8856 15206 8902 15258
rect 8902 15206 8912 15258
rect 8936 15206 8966 15258
rect 8966 15206 8978 15258
rect 8978 15206 8992 15258
rect 9016 15206 9030 15258
rect 9030 15206 9042 15258
rect 9042 15206 9072 15258
rect 9096 15206 9106 15258
rect 9106 15206 9152 15258
rect 8856 15204 8912 15206
rect 8936 15204 8992 15206
rect 9016 15204 9072 15206
rect 9096 15204 9152 15206
rect 5856 13082 5912 13084
rect 5936 13082 5992 13084
rect 6016 13082 6072 13084
rect 6096 13082 6152 13084
rect 5856 13030 5902 13082
rect 5902 13030 5912 13082
rect 5936 13030 5966 13082
rect 5966 13030 5978 13082
rect 5978 13030 5992 13082
rect 6016 13030 6030 13082
rect 6030 13030 6042 13082
rect 6042 13030 6072 13082
rect 6096 13030 6106 13082
rect 6106 13030 6152 13082
rect 5856 13028 5912 13030
rect 5936 13028 5992 13030
rect 6016 13028 6072 13030
rect 6096 13028 6152 13030
rect 6182 12688 6238 12744
rect 5856 11994 5912 11996
rect 5936 11994 5992 11996
rect 6016 11994 6072 11996
rect 6096 11994 6152 11996
rect 5856 11942 5902 11994
rect 5902 11942 5912 11994
rect 5936 11942 5966 11994
rect 5966 11942 5978 11994
rect 5978 11942 5992 11994
rect 6016 11942 6030 11994
rect 6030 11942 6042 11994
rect 6042 11942 6072 11994
rect 6096 11942 6106 11994
rect 6106 11942 6152 11994
rect 5856 11940 5912 11942
rect 5936 11940 5992 11942
rect 6016 11940 6072 11942
rect 6096 11940 6152 11942
rect 5856 10906 5912 10908
rect 5936 10906 5992 10908
rect 6016 10906 6072 10908
rect 6096 10906 6152 10908
rect 5856 10854 5902 10906
rect 5902 10854 5912 10906
rect 5936 10854 5966 10906
rect 5966 10854 5978 10906
rect 5978 10854 5992 10906
rect 6016 10854 6030 10906
rect 6030 10854 6042 10906
rect 6042 10854 6072 10906
rect 6096 10854 6106 10906
rect 6106 10854 6152 10906
rect 5856 10852 5912 10854
rect 5936 10852 5992 10854
rect 6016 10852 6072 10854
rect 6096 10852 6152 10854
rect 8856 14170 8912 14172
rect 8936 14170 8992 14172
rect 9016 14170 9072 14172
rect 9096 14170 9152 14172
rect 8856 14118 8902 14170
rect 8902 14118 8912 14170
rect 8936 14118 8966 14170
rect 8966 14118 8978 14170
rect 8978 14118 8992 14170
rect 9016 14118 9030 14170
rect 9030 14118 9042 14170
rect 9042 14118 9072 14170
rect 9096 14118 9106 14170
rect 9106 14118 9152 14170
rect 8856 14116 8912 14118
rect 8936 14116 8992 14118
rect 9016 14116 9072 14118
rect 9096 14116 9152 14118
rect 10356 14714 10412 14716
rect 10436 14714 10492 14716
rect 10516 14714 10572 14716
rect 10596 14714 10652 14716
rect 10356 14662 10402 14714
rect 10402 14662 10412 14714
rect 10436 14662 10466 14714
rect 10466 14662 10478 14714
rect 10478 14662 10492 14714
rect 10516 14662 10530 14714
rect 10530 14662 10542 14714
rect 10542 14662 10572 14714
rect 10596 14662 10606 14714
rect 10606 14662 10652 14714
rect 10356 14660 10412 14662
rect 10436 14660 10492 14662
rect 10516 14660 10572 14662
rect 10596 14660 10652 14662
rect 8856 13082 8912 13084
rect 8936 13082 8992 13084
rect 9016 13082 9072 13084
rect 9096 13082 9152 13084
rect 8856 13030 8902 13082
rect 8902 13030 8912 13082
rect 8936 13030 8966 13082
rect 8966 13030 8978 13082
rect 8978 13030 8992 13082
rect 9016 13030 9030 13082
rect 9030 13030 9042 13082
rect 9042 13030 9072 13082
rect 9096 13030 9106 13082
rect 9106 13030 9152 13082
rect 8856 13028 8912 13030
rect 8936 13028 8992 13030
rect 9016 13028 9072 13030
rect 9096 13028 9152 13030
rect 6182 10684 6184 10704
rect 6184 10684 6236 10704
rect 6236 10684 6238 10704
rect 6182 10648 6238 10684
rect 5856 9818 5912 9820
rect 5936 9818 5992 9820
rect 6016 9818 6072 9820
rect 6096 9818 6152 9820
rect 5856 9766 5902 9818
rect 5902 9766 5912 9818
rect 5936 9766 5966 9818
rect 5966 9766 5978 9818
rect 5978 9766 5992 9818
rect 6016 9766 6030 9818
rect 6030 9766 6042 9818
rect 6042 9766 6072 9818
rect 6096 9766 6106 9818
rect 6106 9766 6152 9818
rect 5856 9764 5912 9766
rect 5936 9764 5992 9766
rect 6016 9764 6072 9766
rect 6096 9764 6152 9766
rect 7356 12538 7412 12540
rect 7436 12538 7492 12540
rect 7516 12538 7572 12540
rect 7596 12538 7652 12540
rect 7356 12486 7402 12538
rect 7402 12486 7412 12538
rect 7436 12486 7466 12538
rect 7466 12486 7478 12538
rect 7478 12486 7492 12538
rect 7516 12486 7530 12538
rect 7530 12486 7542 12538
rect 7542 12486 7572 12538
rect 7596 12486 7606 12538
rect 7606 12486 7652 12538
rect 7356 12484 7412 12486
rect 7436 12484 7492 12486
rect 7516 12484 7572 12486
rect 7596 12484 7652 12486
rect 7356 11450 7412 11452
rect 7436 11450 7492 11452
rect 7516 11450 7572 11452
rect 7596 11450 7652 11452
rect 7356 11398 7402 11450
rect 7402 11398 7412 11450
rect 7436 11398 7466 11450
rect 7466 11398 7478 11450
rect 7478 11398 7492 11450
rect 7516 11398 7530 11450
rect 7530 11398 7542 11450
rect 7542 11398 7572 11450
rect 7596 11398 7606 11450
rect 7606 11398 7652 11450
rect 7356 11396 7412 11398
rect 7436 11396 7492 11398
rect 7516 11396 7572 11398
rect 7596 11396 7652 11398
rect 8206 10648 8262 10704
rect 7356 10362 7412 10364
rect 7436 10362 7492 10364
rect 7516 10362 7572 10364
rect 7596 10362 7652 10364
rect 7356 10310 7402 10362
rect 7402 10310 7412 10362
rect 7436 10310 7466 10362
rect 7466 10310 7478 10362
rect 7478 10310 7492 10362
rect 7516 10310 7530 10362
rect 7530 10310 7542 10362
rect 7542 10310 7572 10362
rect 7596 10310 7606 10362
rect 7606 10310 7652 10362
rect 7356 10308 7412 10310
rect 7436 10308 7492 10310
rect 7516 10308 7572 10310
rect 7596 10308 7652 10310
rect 8856 11994 8912 11996
rect 8936 11994 8992 11996
rect 9016 11994 9072 11996
rect 9096 11994 9152 11996
rect 8856 11942 8902 11994
rect 8902 11942 8912 11994
rect 8936 11942 8966 11994
rect 8966 11942 8978 11994
rect 8978 11942 8992 11994
rect 9016 11942 9030 11994
rect 9030 11942 9042 11994
rect 9042 11942 9072 11994
rect 9096 11942 9106 11994
rect 9106 11942 9152 11994
rect 8856 11940 8912 11942
rect 8936 11940 8992 11942
rect 9016 11940 9072 11942
rect 9096 11940 9152 11942
rect 8942 11076 8998 11112
rect 8942 11056 8944 11076
rect 8944 11056 8996 11076
rect 8996 11056 8998 11076
rect 8856 10906 8912 10908
rect 8936 10906 8992 10908
rect 9016 10906 9072 10908
rect 9096 10906 9152 10908
rect 8856 10854 8902 10906
rect 8902 10854 8912 10906
rect 8936 10854 8966 10906
rect 8966 10854 8978 10906
rect 8978 10854 8992 10906
rect 9016 10854 9030 10906
rect 9030 10854 9042 10906
rect 9042 10854 9072 10906
rect 9096 10854 9106 10906
rect 9106 10854 9152 10906
rect 8856 10852 8912 10854
rect 8936 10852 8992 10854
rect 9016 10852 9072 10854
rect 9096 10852 9152 10854
rect 11856 23962 11912 23964
rect 11936 23962 11992 23964
rect 12016 23962 12072 23964
rect 12096 23962 12152 23964
rect 11856 23910 11902 23962
rect 11902 23910 11912 23962
rect 11936 23910 11966 23962
rect 11966 23910 11978 23962
rect 11978 23910 11992 23962
rect 12016 23910 12030 23962
rect 12030 23910 12042 23962
rect 12042 23910 12072 23962
rect 12096 23910 12106 23962
rect 12106 23910 12152 23962
rect 11856 23908 11912 23910
rect 11936 23908 11992 23910
rect 12016 23908 12072 23910
rect 12096 23908 12152 23910
rect 11856 22874 11912 22876
rect 11936 22874 11992 22876
rect 12016 22874 12072 22876
rect 12096 22874 12152 22876
rect 11856 22822 11902 22874
rect 11902 22822 11912 22874
rect 11936 22822 11966 22874
rect 11966 22822 11978 22874
rect 11978 22822 11992 22874
rect 12016 22822 12030 22874
rect 12030 22822 12042 22874
rect 12042 22822 12072 22874
rect 12096 22822 12106 22874
rect 12106 22822 12152 22874
rect 11856 22820 11912 22822
rect 11936 22820 11992 22822
rect 12016 22820 12072 22822
rect 12096 22820 12152 22822
rect 11856 21786 11912 21788
rect 11936 21786 11992 21788
rect 12016 21786 12072 21788
rect 12096 21786 12152 21788
rect 11856 21734 11902 21786
rect 11902 21734 11912 21786
rect 11936 21734 11966 21786
rect 11966 21734 11978 21786
rect 11978 21734 11992 21786
rect 12016 21734 12030 21786
rect 12030 21734 12042 21786
rect 12042 21734 12072 21786
rect 12096 21734 12106 21786
rect 12106 21734 12152 21786
rect 11856 21732 11912 21734
rect 11936 21732 11992 21734
rect 12016 21732 12072 21734
rect 12096 21732 12152 21734
rect 11856 20698 11912 20700
rect 11936 20698 11992 20700
rect 12016 20698 12072 20700
rect 12096 20698 12152 20700
rect 11856 20646 11902 20698
rect 11902 20646 11912 20698
rect 11936 20646 11966 20698
rect 11966 20646 11978 20698
rect 11978 20646 11992 20698
rect 12016 20646 12030 20698
rect 12030 20646 12042 20698
rect 12042 20646 12072 20698
rect 12096 20646 12106 20698
rect 12106 20646 12152 20698
rect 11856 20644 11912 20646
rect 11936 20644 11992 20646
rect 12016 20644 12072 20646
rect 12096 20644 12152 20646
rect 11856 19610 11912 19612
rect 11936 19610 11992 19612
rect 12016 19610 12072 19612
rect 12096 19610 12152 19612
rect 11856 19558 11902 19610
rect 11902 19558 11912 19610
rect 11936 19558 11966 19610
rect 11966 19558 11978 19610
rect 11978 19558 11992 19610
rect 12016 19558 12030 19610
rect 12030 19558 12042 19610
rect 12042 19558 12072 19610
rect 12096 19558 12106 19610
rect 12106 19558 12152 19610
rect 11856 19556 11912 19558
rect 11936 19556 11992 19558
rect 12016 19556 12072 19558
rect 12096 19556 12152 19558
rect 11856 18522 11912 18524
rect 11936 18522 11992 18524
rect 12016 18522 12072 18524
rect 12096 18522 12152 18524
rect 11856 18470 11902 18522
rect 11902 18470 11912 18522
rect 11936 18470 11966 18522
rect 11966 18470 11978 18522
rect 11978 18470 11992 18522
rect 12016 18470 12030 18522
rect 12030 18470 12042 18522
rect 12042 18470 12072 18522
rect 12096 18470 12106 18522
rect 12106 18470 12152 18522
rect 11856 18468 11912 18470
rect 11936 18468 11992 18470
rect 12016 18468 12072 18470
rect 12096 18468 12152 18470
rect 11856 17434 11912 17436
rect 11936 17434 11992 17436
rect 12016 17434 12072 17436
rect 12096 17434 12152 17436
rect 11856 17382 11902 17434
rect 11902 17382 11912 17434
rect 11936 17382 11966 17434
rect 11966 17382 11978 17434
rect 11978 17382 11992 17434
rect 12016 17382 12030 17434
rect 12030 17382 12042 17434
rect 12042 17382 12072 17434
rect 12096 17382 12106 17434
rect 12106 17382 12152 17434
rect 11856 17380 11912 17382
rect 11936 17380 11992 17382
rect 12016 17380 12072 17382
rect 12096 17380 12152 17382
rect 11856 16346 11912 16348
rect 11936 16346 11992 16348
rect 12016 16346 12072 16348
rect 12096 16346 12152 16348
rect 11856 16294 11902 16346
rect 11902 16294 11912 16346
rect 11936 16294 11966 16346
rect 11966 16294 11978 16346
rect 11978 16294 11992 16346
rect 12016 16294 12030 16346
rect 12030 16294 12042 16346
rect 12042 16294 12072 16346
rect 12096 16294 12106 16346
rect 12106 16294 12152 16346
rect 11856 16292 11912 16294
rect 11936 16292 11992 16294
rect 12016 16292 12072 16294
rect 12096 16292 12152 16294
rect 10356 13626 10412 13628
rect 10436 13626 10492 13628
rect 10516 13626 10572 13628
rect 10596 13626 10652 13628
rect 10356 13574 10402 13626
rect 10402 13574 10412 13626
rect 10436 13574 10466 13626
rect 10466 13574 10478 13626
rect 10478 13574 10492 13626
rect 10516 13574 10530 13626
rect 10530 13574 10542 13626
rect 10542 13574 10572 13626
rect 10596 13574 10606 13626
rect 10606 13574 10652 13626
rect 10356 13572 10412 13574
rect 10436 13572 10492 13574
rect 10516 13572 10572 13574
rect 10596 13572 10652 13574
rect 10356 12538 10412 12540
rect 10436 12538 10492 12540
rect 10516 12538 10572 12540
rect 10596 12538 10652 12540
rect 10356 12486 10402 12538
rect 10402 12486 10412 12538
rect 10436 12486 10466 12538
rect 10466 12486 10478 12538
rect 10478 12486 10492 12538
rect 10516 12486 10530 12538
rect 10530 12486 10542 12538
rect 10542 12486 10572 12538
rect 10596 12486 10606 12538
rect 10606 12486 10652 12538
rect 10356 12484 10412 12486
rect 10436 12484 10492 12486
rect 10516 12484 10572 12486
rect 10596 12484 10652 12486
rect 11856 15258 11912 15260
rect 11936 15258 11992 15260
rect 12016 15258 12072 15260
rect 12096 15258 12152 15260
rect 11856 15206 11902 15258
rect 11902 15206 11912 15258
rect 11936 15206 11966 15258
rect 11966 15206 11978 15258
rect 11978 15206 11992 15258
rect 12016 15206 12030 15258
rect 12030 15206 12042 15258
rect 12042 15206 12072 15258
rect 12096 15206 12106 15258
rect 12106 15206 12152 15258
rect 11856 15204 11912 15206
rect 11936 15204 11992 15206
rect 12016 15204 12072 15206
rect 12096 15204 12152 15206
rect 11856 14170 11912 14172
rect 11936 14170 11992 14172
rect 12016 14170 12072 14172
rect 12096 14170 12152 14172
rect 11856 14118 11902 14170
rect 11902 14118 11912 14170
rect 11936 14118 11966 14170
rect 11966 14118 11978 14170
rect 11978 14118 11992 14170
rect 12016 14118 12030 14170
rect 12030 14118 12042 14170
rect 12042 14118 12072 14170
rect 12096 14118 12106 14170
rect 12106 14118 12152 14170
rect 11856 14116 11912 14118
rect 11936 14116 11992 14118
rect 12016 14116 12072 14118
rect 12096 14116 12152 14118
rect 12530 13948 12532 13968
rect 12532 13948 12584 13968
rect 12584 13948 12586 13968
rect 12530 13912 12586 13948
rect 10356 11450 10412 11452
rect 10436 11450 10492 11452
rect 10516 11450 10572 11452
rect 10596 11450 10652 11452
rect 10356 11398 10402 11450
rect 10402 11398 10412 11450
rect 10436 11398 10466 11450
rect 10466 11398 10478 11450
rect 10478 11398 10492 11450
rect 10516 11398 10530 11450
rect 10530 11398 10542 11450
rect 10542 11398 10572 11450
rect 10596 11398 10606 11450
rect 10606 11398 10652 11450
rect 10356 11396 10412 11398
rect 10436 11396 10492 11398
rect 10516 11396 10572 11398
rect 10596 11396 10652 11398
rect 7356 9274 7412 9276
rect 7436 9274 7492 9276
rect 7516 9274 7572 9276
rect 7596 9274 7652 9276
rect 7356 9222 7402 9274
rect 7402 9222 7412 9274
rect 7436 9222 7466 9274
rect 7466 9222 7478 9274
rect 7478 9222 7492 9274
rect 7516 9222 7530 9274
rect 7530 9222 7542 9274
rect 7542 9222 7572 9274
rect 7596 9222 7606 9274
rect 7606 9222 7652 9274
rect 7356 9220 7412 9222
rect 7436 9220 7492 9222
rect 7516 9220 7572 9222
rect 7596 9220 7652 9222
rect 8856 9818 8912 9820
rect 8936 9818 8992 9820
rect 9016 9818 9072 9820
rect 9096 9818 9152 9820
rect 8856 9766 8902 9818
rect 8902 9766 8912 9818
rect 8936 9766 8966 9818
rect 8966 9766 8978 9818
rect 8978 9766 8992 9818
rect 9016 9766 9030 9818
rect 9030 9766 9042 9818
rect 9042 9766 9072 9818
rect 9096 9766 9106 9818
rect 9106 9766 9152 9818
rect 8856 9764 8912 9766
rect 8936 9764 8992 9766
rect 9016 9764 9072 9766
rect 9096 9764 9152 9766
rect 10356 10362 10412 10364
rect 10436 10362 10492 10364
rect 10516 10362 10572 10364
rect 10596 10362 10652 10364
rect 10356 10310 10402 10362
rect 10402 10310 10412 10362
rect 10436 10310 10466 10362
rect 10466 10310 10478 10362
rect 10478 10310 10492 10362
rect 10516 10310 10530 10362
rect 10530 10310 10542 10362
rect 10542 10310 10572 10362
rect 10596 10310 10606 10362
rect 10606 10310 10652 10362
rect 10356 10308 10412 10310
rect 10436 10308 10492 10310
rect 10516 10308 10572 10310
rect 10596 10308 10652 10310
rect 4356 8186 4412 8188
rect 4436 8186 4492 8188
rect 4516 8186 4572 8188
rect 4596 8186 4652 8188
rect 4356 8134 4402 8186
rect 4402 8134 4412 8186
rect 4436 8134 4466 8186
rect 4466 8134 4478 8186
rect 4478 8134 4492 8186
rect 4516 8134 4530 8186
rect 4530 8134 4542 8186
rect 4542 8134 4572 8186
rect 4596 8134 4606 8186
rect 4606 8134 4652 8186
rect 4356 8132 4412 8134
rect 4436 8132 4492 8134
rect 4516 8132 4572 8134
rect 4596 8132 4652 8134
rect 1356 7098 1412 7100
rect 1436 7098 1492 7100
rect 1516 7098 1572 7100
rect 1596 7098 1652 7100
rect 1356 7046 1402 7098
rect 1402 7046 1412 7098
rect 1436 7046 1466 7098
rect 1466 7046 1478 7098
rect 1478 7046 1492 7098
rect 1516 7046 1530 7098
rect 1530 7046 1542 7098
rect 1542 7046 1572 7098
rect 1596 7046 1606 7098
rect 1606 7046 1652 7098
rect 1356 7044 1412 7046
rect 1436 7044 1492 7046
rect 1516 7044 1572 7046
rect 1596 7044 1652 7046
rect 5856 8730 5912 8732
rect 5936 8730 5992 8732
rect 6016 8730 6072 8732
rect 6096 8730 6152 8732
rect 5856 8678 5902 8730
rect 5902 8678 5912 8730
rect 5936 8678 5966 8730
rect 5966 8678 5978 8730
rect 5978 8678 5992 8730
rect 6016 8678 6030 8730
rect 6030 8678 6042 8730
rect 6042 8678 6072 8730
rect 6096 8678 6106 8730
rect 6106 8678 6152 8730
rect 5856 8676 5912 8678
rect 5936 8676 5992 8678
rect 6016 8676 6072 8678
rect 6096 8676 6152 8678
rect 7356 8186 7412 8188
rect 7436 8186 7492 8188
rect 7516 8186 7572 8188
rect 7596 8186 7652 8188
rect 7356 8134 7402 8186
rect 7402 8134 7412 8186
rect 7436 8134 7466 8186
rect 7466 8134 7478 8186
rect 7478 8134 7492 8186
rect 7516 8134 7530 8186
rect 7530 8134 7542 8186
rect 7542 8134 7572 8186
rect 7596 8134 7606 8186
rect 7606 8134 7652 8186
rect 7356 8132 7412 8134
rect 7436 8132 7492 8134
rect 7516 8132 7572 8134
rect 7596 8132 7652 8134
rect 5856 7642 5912 7644
rect 5936 7642 5992 7644
rect 6016 7642 6072 7644
rect 6096 7642 6152 7644
rect 5856 7590 5902 7642
rect 5902 7590 5912 7642
rect 5936 7590 5966 7642
rect 5966 7590 5978 7642
rect 5978 7590 5992 7642
rect 6016 7590 6030 7642
rect 6030 7590 6042 7642
rect 6042 7590 6072 7642
rect 6096 7590 6106 7642
rect 6106 7590 6152 7642
rect 5856 7588 5912 7590
rect 5936 7588 5992 7590
rect 6016 7588 6072 7590
rect 6096 7588 6152 7590
rect 4356 7098 4412 7100
rect 4436 7098 4492 7100
rect 4516 7098 4572 7100
rect 4596 7098 4652 7100
rect 4356 7046 4402 7098
rect 4402 7046 4412 7098
rect 4436 7046 4466 7098
rect 4466 7046 4478 7098
rect 4478 7046 4492 7098
rect 4516 7046 4530 7098
rect 4530 7046 4542 7098
rect 4542 7046 4572 7098
rect 4596 7046 4606 7098
rect 4606 7046 4652 7098
rect 4356 7044 4412 7046
rect 4436 7044 4492 7046
rect 4516 7044 4572 7046
rect 4596 7044 4652 7046
rect 2856 6554 2912 6556
rect 2936 6554 2992 6556
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 2856 6502 2902 6554
rect 2902 6502 2912 6554
rect 2936 6502 2966 6554
rect 2966 6502 2978 6554
rect 2978 6502 2992 6554
rect 3016 6502 3030 6554
rect 3030 6502 3042 6554
rect 3042 6502 3072 6554
rect 3096 6502 3106 6554
rect 3106 6502 3152 6554
rect 2856 6500 2912 6502
rect 2936 6500 2992 6502
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 1356 6010 1412 6012
rect 1436 6010 1492 6012
rect 1516 6010 1572 6012
rect 1596 6010 1652 6012
rect 1356 5958 1402 6010
rect 1402 5958 1412 6010
rect 1436 5958 1466 6010
rect 1466 5958 1478 6010
rect 1478 5958 1492 6010
rect 1516 5958 1530 6010
rect 1530 5958 1542 6010
rect 1542 5958 1572 6010
rect 1596 5958 1606 6010
rect 1606 5958 1652 6010
rect 1356 5956 1412 5958
rect 1436 5956 1492 5958
rect 1516 5956 1572 5958
rect 1596 5956 1652 5958
rect 4356 6010 4412 6012
rect 4436 6010 4492 6012
rect 4516 6010 4572 6012
rect 4596 6010 4652 6012
rect 4356 5958 4402 6010
rect 4402 5958 4412 6010
rect 4436 5958 4466 6010
rect 4466 5958 4478 6010
rect 4478 5958 4492 6010
rect 4516 5958 4530 6010
rect 4530 5958 4542 6010
rect 4542 5958 4572 6010
rect 4596 5958 4606 6010
rect 4606 5958 4652 6010
rect 4356 5956 4412 5958
rect 4436 5956 4492 5958
rect 4516 5956 4572 5958
rect 4596 5956 4652 5958
rect 5856 6554 5912 6556
rect 5936 6554 5992 6556
rect 6016 6554 6072 6556
rect 6096 6554 6152 6556
rect 5856 6502 5902 6554
rect 5902 6502 5912 6554
rect 5936 6502 5966 6554
rect 5966 6502 5978 6554
rect 5978 6502 5992 6554
rect 6016 6502 6030 6554
rect 6030 6502 6042 6554
rect 6042 6502 6072 6554
rect 6096 6502 6106 6554
rect 6106 6502 6152 6554
rect 5856 6500 5912 6502
rect 5936 6500 5992 6502
rect 6016 6500 6072 6502
rect 6096 6500 6152 6502
rect 2856 5466 2912 5468
rect 2936 5466 2992 5468
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 2856 5414 2902 5466
rect 2902 5414 2912 5466
rect 2936 5414 2966 5466
rect 2966 5414 2978 5466
rect 2978 5414 2992 5466
rect 3016 5414 3030 5466
rect 3030 5414 3042 5466
rect 3042 5414 3072 5466
rect 3096 5414 3106 5466
rect 3106 5414 3152 5466
rect 2856 5412 2912 5414
rect 2936 5412 2992 5414
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 1356 4922 1412 4924
rect 1436 4922 1492 4924
rect 1516 4922 1572 4924
rect 1596 4922 1652 4924
rect 1356 4870 1402 4922
rect 1402 4870 1412 4922
rect 1436 4870 1466 4922
rect 1466 4870 1478 4922
rect 1478 4870 1492 4922
rect 1516 4870 1530 4922
rect 1530 4870 1542 4922
rect 1542 4870 1572 4922
rect 1596 4870 1606 4922
rect 1606 4870 1652 4922
rect 1356 4868 1412 4870
rect 1436 4868 1492 4870
rect 1516 4868 1572 4870
rect 1596 4868 1652 4870
rect 4356 4922 4412 4924
rect 4436 4922 4492 4924
rect 4516 4922 4572 4924
rect 4596 4922 4652 4924
rect 4356 4870 4402 4922
rect 4402 4870 4412 4922
rect 4436 4870 4466 4922
rect 4466 4870 4478 4922
rect 4478 4870 4492 4922
rect 4516 4870 4530 4922
rect 4530 4870 4542 4922
rect 4542 4870 4572 4922
rect 4596 4870 4606 4922
rect 4606 4870 4652 4922
rect 4356 4868 4412 4870
rect 4436 4868 4492 4870
rect 4516 4868 4572 4870
rect 4596 4868 4652 4870
rect 2856 4378 2912 4380
rect 2936 4378 2992 4380
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 2856 4326 2902 4378
rect 2902 4326 2912 4378
rect 2936 4326 2966 4378
rect 2966 4326 2978 4378
rect 2978 4326 2992 4378
rect 3016 4326 3030 4378
rect 3030 4326 3042 4378
rect 3042 4326 3072 4378
rect 3096 4326 3106 4378
rect 3106 4326 3152 4378
rect 2856 4324 2912 4326
rect 2936 4324 2992 4326
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 1356 3834 1412 3836
rect 1436 3834 1492 3836
rect 1516 3834 1572 3836
rect 1596 3834 1652 3836
rect 1356 3782 1402 3834
rect 1402 3782 1412 3834
rect 1436 3782 1466 3834
rect 1466 3782 1478 3834
rect 1478 3782 1492 3834
rect 1516 3782 1530 3834
rect 1530 3782 1542 3834
rect 1542 3782 1572 3834
rect 1596 3782 1606 3834
rect 1606 3782 1652 3834
rect 1356 3780 1412 3782
rect 1436 3780 1492 3782
rect 1516 3780 1572 3782
rect 1596 3780 1652 3782
rect 4356 3834 4412 3836
rect 4436 3834 4492 3836
rect 4516 3834 4572 3836
rect 4596 3834 4652 3836
rect 4356 3782 4402 3834
rect 4402 3782 4412 3834
rect 4436 3782 4466 3834
rect 4466 3782 4478 3834
rect 4478 3782 4492 3834
rect 4516 3782 4530 3834
rect 4530 3782 4542 3834
rect 4542 3782 4572 3834
rect 4596 3782 4606 3834
rect 4606 3782 4652 3834
rect 4356 3780 4412 3782
rect 4436 3780 4492 3782
rect 4516 3780 4572 3782
rect 4596 3780 4652 3782
rect 5856 5466 5912 5468
rect 5936 5466 5992 5468
rect 6016 5466 6072 5468
rect 6096 5466 6152 5468
rect 5856 5414 5902 5466
rect 5902 5414 5912 5466
rect 5936 5414 5966 5466
rect 5966 5414 5978 5466
rect 5978 5414 5992 5466
rect 6016 5414 6030 5466
rect 6030 5414 6042 5466
rect 6042 5414 6072 5466
rect 6096 5414 6106 5466
rect 6106 5414 6152 5466
rect 5856 5412 5912 5414
rect 5936 5412 5992 5414
rect 6016 5412 6072 5414
rect 6096 5412 6152 5414
rect 5856 4378 5912 4380
rect 5936 4378 5992 4380
rect 6016 4378 6072 4380
rect 6096 4378 6152 4380
rect 5856 4326 5902 4378
rect 5902 4326 5912 4378
rect 5936 4326 5966 4378
rect 5966 4326 5978 4378
rect 5978 4326 5992 4378
rect 6016 4326 6030 4378
rect 6030 4326 6042 4378
rect 6042 4326 6072 4378
rect 6096 4326 6106 4378
rect 6106 4326 6152 4378
rect 5856 4324 5912 4326
rect 5936 4324 5992 4326
rect 6016 4324 6072 4326
rect 6096 4324 6152 4326
rect 2856 3290 2912 3292
rect 2936 3290 2992 3292
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 2856 3238 2902 3290
rect 2902 3238 2912 3290
rect 2936 3238 2966 3290
rect 2966 3238 2978 3290
rect 2978 3238 2992 3290
rect 3016 3238 3030 3290
rect 3030 3238 3042 3290
rect 3042 3238 3072 3290
rect 3096 3238 3106 3290
rect 3106 3238 3152 3290
rect 2856 3236 2912 3238
rect 2936 3236 2992 3238
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 5856 3290 5912 3292
rect 5936 3290 5992 3292
rect 6016 3290 6072 3292
rect 6096 3290 6152 3292
rect 5856 3238 5902 3290
rect 5902 3238 5912 3290
rect 5936 3238 5966 3290
rect 5966 3238 5978 3290
rect 5978 3238 5992 3290
rect 6016 3238 6030 3290
rect 6030 3238 6042 3290
rect 6042 3238 6072 3290
rect 6096 3238 6106 3290
rect 6106 3238 6152 3290
rect 5856 3236 5912 3238
rect 5936 3236 5992 3238
rect 6016 3236 6072 3238
rect 6096 3236 6152 3238
rect 7356 7098 7412 7100
rect 7436 7098 7492 7100
rect 7516 7098 7572 7100
rect 7596 7098 7652 7100
rect 7356 7046 7402 7098
rect 7402 7046 7412 7098
rect 7436 7046 7466 7098
rect 7466 7046 7478 7098
rect 7478 7046 7492 7098
rect 7516 7046 7530 7098
rect 7530 7046 7542 7098
rect 7542 7046 7572 7098
rect 7596 7046 7606 7098
rect 7606 7046 7652 7098
rect 7356 7044 7412 7046
rect 7436 7044 7492 7046
rect 7516 7044 7572 7046
rect 7596 7044 7652 7046
rect 7356 6010 7412 6012
rect 7436 6010 7492 6012
rect 7516 6010 7572 6012
rect 7596 6010 7652 6012
rect 7356 5958 7402 6010
rect 7402 5958 7412 6010
rect 7436 5958 7466 6010
rect 7466 5958 7478 6010
rect 7478 5958 7492 6010
rect 7516 5958 7530 6010
rect 7530 5958 7542 6010
rect 7542 5958 7572 6010
rect 7596 5958 7606 6010
rect 7606 5958 7652 6010
rect 7356 5956 7412 5958
rect 7436 5956 7492 5958
rect 7516 5956 7572 5958
rect 7596 5956 7652 5958
rect 1356 2746 1412 2748
rect 1436 2746 1492 2748
rect 1516 2746 1572 2748
rect 1596 2746 1652 2748
rect 1356 2694 1402 2746
rect 1402 2694 1412 2746
rect 1436 2694 1466 2746
rect 1466 2694 1478 2746
rect 1478 2694 1492 2746
rect 1516 2694 1530 2746
rect 1530 2694 1542 2746
rect 1542 2694 1572 2746
rect 1596 2694 1606 2746
rect 1606 2694 1652 2746
rect 1356 2692 1412 2694
rect 1436 2692 1492 2694
rect 1516 2692 1572 2694
rect 1596 2692 1652 2694
rect 4356 2746 4412 2748
rect 4436 2746 4492 2748
rect 4516 2746 4572 2748
rect 4596 2746 4652 2748
rect 4356 2694 4402 2746
rect 4402 2694 4412 2746
rect 4436 2694 4466 2746
rect 4466 2694 4478 2746
rect 4478 2694 4492 2746
rect 4516 2694 4530 2746
rect 4530 2694 4542 2746
rect 4542 2694 4572 2746
rect 4596 2694 4606 2746
rect 4606 2694 4652 2746
rect 4356 2692 4412 2694
rect 4436 2692 4492 2694
rect 4516 2692 4572 2694
rect 4596 2692 4652 2694
rect 8856 8730 8912 8732
rect 8936 8730 8992 8732
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 8856 8678 8902 8730
rect 8902 8678 8912 8730
rect 8936 8678 8966 8730
rect 8966 8678 8978 8730
rect 8978 8678 8992 8730
rect 9016 8678 9030 8730
rect 9030 8678 9042 8730
rect 9042 8678 9072 8730
rect 9096 8678 9106 8730
rect 9106 8678 9152 8730
rect 8856 8676 8912 8678
rect 8936 8676 8992 8678
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 8856 7642 8912 7644
rect 8936 7642 8992 7644
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 8856 7590 8902 7642
rect 8902 7590 8912 7642
rect 8936 7590 8966 7642
rect 8966 7590 8978 7642
rect 8978 7590 8992 7642
rect 9016 7590 9030 7642
rect 9030 7590 9042 7642
rect 9042 7590 9072 7642
rect 9096 7590 9106 7642
rect 9106 7590 9152 7642
rect 8856 7588 8912 7590
rect 8936 7588 8992 7590
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 7356 4922 7412 4924
rect 7436 4922 7492 4924
rect 7516 4922 7572 4924
rect 7596 4922 7652 4924
rect 7356 4870 7402 4922
rect 7402 4870 7412 4922
rect 7436 4870 7466 4922
rect 7466 4870 7478 4922
rect 7478 4870 7492 4922
rect 7516 4870 7530 4922
rect 7530 4870 7542 4922
rect 7542 4870 7572 4922
rect 7596 4870 7606 4922
rect 7606 4870 7652 4922
rect 7356 4868 7412 4870
rect 7436 4868 7492 4870
rect 7516 4868 7572 4870
rect 7596 4868 7652 4870
rect 7356 3834 7412 3836
rect 7436 3834 7492 3836
rect 7516 3834 7572 3836
rect 7596 3834 7652 3836
rect 7356 3782 7402 3834
rect 7402 3782 7412 3834
rect 7436 3782 7466 3834
rect 7466 3782 7478 3834
rect 7478 3782 7492 3834
rect 7516 3782 7530 3834
rect 7530 3782 7542 3834
rect 7542 3782 7572 3834
rect 7596 3782 7606 3834
rect 7606 3782 7652 3834
rect 7356 3780 7412 3782
rect 7436 3780 7492 3782
rect 7516 3780 7572 3782
rect 7596 3780 7652 3782
rect 7356 2746 7412 2748
rect 7436 2746 7492 2748
rect 7516 2746 7572 2748
rect 7596 2746 7652 2748
rect 7356 2694 7402 2746
rect 7402 2694 7412 2746
rect 7436 2694 7466 2746
rect 7466 2694 7478 2746
rect 7478 2694 7492 2746
rect 7516 2694 7530 2746
rect 7530 2694 7542 2746
rect 7542 2694 7572 2746
rect 7596 2694 7606 2746
rect 7606 2694 7652 2746
rect 7356 2692 7412 2694
rect 7436 2692 7492 2694
rect 7516 2692 7572 2694
rect 7596 2692 7652 2694
rect 8856 6554 8912 6556
rect 8936 6554 8992 6556
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 8856 6502 8902 6554
rect 8902 6502 8912 6554
rect 8936 6502 8966 6554
rect 8966 6502 8978 6554
rect 8978 6502 8992 6554
rect 9016 6502 9030 6554
rect 9030 6502 9042 6554
rect 9042 6502 9072 6554
rect 9096 6502 9106 6554
rect 9106 6502 9152 6554
rect 8856 6500 8912 6502
rect 8936 6500 8992 6502
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 10356 9274 10412 9276
rect 10436 9274 10492 9276
rect 10516 9274 10572 9276
rect 10596 9274 10652 9276
rect 10356 9222 10402 9274
rect 10402 9222 10412 9274
rect 10436 9222 10466 9274
rect 10466 9222 10478 9274
rect 10478 9222 10492 9274
rect 10516 9222 10530 9274
rect 10530 9222 10542 9274
rect 10542 9222 10572 9274
rect 10596 9222 10606 9274
rect 10606 9222 10652 9274
rect 10356 9220 10412 9222
rect 10436 9220 10492 9222
rect 10516 9220 10572 9222
rect 10596 9220 10652 9222
rect 10356 8186 10412 8188
rect 10436 8186 10492 8188
rect 10516 8186 10572 8188
rect 10596 8186 10652 8188
rect 10356 8134 10402 8186
rect 10402 8134 10412 8186
rect 10436 8134 10466 8186
rect 10466 8134 10478 8186
rect 10478 8134 10492 8186
rect 10516 8134 10530 8186
rect 10530 8134 10542 8186
rect 10542 8134 10572 8186
rect 10596 8134 10606 8186
rect 10606 8134 10652 8186
rect 10356 8132 10412 8134
rect 10436 8132 10492 8134
rect 10516 8132 10572 8134
rect 10596 8132 10652 8134
rect 10356 7098 10412 7100
rect 10436 7098 10492 7100
rect 10516 7098 10572 7100
rect 10596 7098 10652 7100
rect 10356 7046 10402 7098
rect 10402 7046 10412 7098
rect 10436 7046 10466 7098
rect 10466 7046 10478 7098
rect 10478 7046 10492 7098
rect 10516 7046 10530 7098
rect 10530 7046 10542 7098
rect 10542 7046 10572 7098
rect 10596 7046 10606 7098
rect 10606 7046 10652 7098
rect 10356 7044 10412 7046
rect 10436 7044 10492 7046
rect 10516 7044 10572 7046
rect 10596 7044 10652 7046
rect 11856 13082 11912 13084
rect 11936 13082 11992 13084
rect 12016 13082 12072 13084
rect 12096 13082 12152 13084
rect 11856 13030 11902 13082
rect 11902 13030 11912 13082
rect 11936 13030 11966 13082
rect 11966 13030 11978 13082
rect 11978 13030 11992 13082
rect 12016 13030 12030 13082
rect 12030 13030 12042 13082
rect 12042 13030 12072 13082
rect 12096 13030 12106 13082
rect 12106 13030 12152 13082
rect 11856 13028 11912 13030
rect 11936 13028 11992 13030
rect 12016 13028 12072 13030
rect 12096 13028 12152 13030
rect 13356 24506 13412 24508
rect 13436 24506 13492 24508
rect 13516 24506 13572 24508
rect 13596 24506 13652 24508
rect 13356 24454 13402 24506
rect 13402 24454 13412 24506
rect 13436 24454 13466 24506
rect 13466 24454 13478 24506
rect 13478 24454 13492 24506
rect 13516 24454 13530 24506
rect 13530 24454 13542 24506
rect 13542 24454 13572 24506
rect 13596 24454 13606 24506
rect 13606 24454 13652 24506
rect 13356 24452 13412 24454
rect 13436 24452 13492 24454
rect 13516 24452 13572 24454
rect 13596 24452 13652 24454
rect 13356 23418 13412 23420
rect 13436 23418 13492 23420
rect 13516 23418 13572 23420
rect 13596 23418 13652 23420
rect 13356 23366 13402 23418
rect 13402 23366 13412 23418
rect 13436 23366 13466 23418
rect 13466 23366 13478 23418
rect 13478 23366 13492 23418
rect 13516 23366 13530 23418
rect 13530 23366 13542 23418
rect 13542 23366 13572 23418
rect 13596 23366 13606 23418
rect 13606 23366 13652 23418
rect 13356 23364 13412 23366
rect 13436 23364 13492 23366
rect 13516 23364 13572 23366
rect 13596 23364 13652 23366
rect 13356 22330 13412 22332
rect 13436 22330 13492 22332
rect 13516 22330 13572 22332
rect 13596 22330 13652 22332
rect 13356 22278 13402 22330
rect 13402 22278 13412 22330
rect 13436 22278 13466 22330
rect 13466 22278 13478 22330
rect 13478 22278 13492 22330
rect 13516 22278 13530 22330
rect 13530 22278 13542 22330
rect 13542 22278 13572 22330
rect 13596 22278 13606 22330
rect 13606 22278 13652 22330
rect 13356 22276 13412 22278
rect 13436 22276 13492 22278
rect 13516 22276 13572 22278
rect 13596 22276 13652 22278
rect 14856 25050 14912 25052
rect 14936 25050 14992 25052
rect 15016 25050 15072 25052
rect 15096 25050 15152 25052
rect 14856 24998 14902 25050
rect 14902 24998 14912 25050
rect 14936 24998 14966 25050
rect 14966 24998 14978 25050
rect 14978 24998 14992 25050
rect 15016 24998 15030 25050
rect 15030 24998 15042 25050
rect 15042 24998 15072 25050
rect 15096 24998 15106 25050
rect 15106 24998 15152 25050
rect 14856 24996 14912 24998
rect 14936 24996 14992 24998
rect 15016 24996 15072 24998
rect 15096 24996 15152 24998
rect 14094 23568 14150 23624
rect 13356 21242 13412 21244
rect 13436 21242 13492 21244
rect 13516 21242 13572 21244
rect 13596 21242 13652 21244
rect 13356 21190 13402 21242
rect 13402 21190 13412 21242
rect 13436 21190 13466 21242
rect 13466 21190 13478 21242
rect 13478 21190 13492 21242
rect 13516 21190 13530 21242
rect 13530 21190 13542 21242
rect 13542 21190 13572 21242
rect 13596 21190 13606 21242
rect 13606 21190 13652 21242
rect 13356 21188 13412 21190
rect 13436 21188 13492 21190
rect 13516 21188 13572 21190
rect 13596 21188 13652 21190
rect 13634 21020 13636 21040
rect 13636 21020 13688 21040
rect 13688 21020 13690 21040
rect 13634 20984 13690 21020
rect 13356 20154 13412 20156
rect 13436 20154 13492 20156
rect 13516 20154 13572 20156
rect 13596 20154 13652 20156
rect 13356 20102 13402 20154
rect 13402 20102 13412 20154
rect 13436 20102 13466 20154
rect 13466 20102 13478 20154
rect 13478 20102 13492 20154
rect 13516 20102 13530 20154
rect 13530 20102 13542 20154
rect 13542 20102 13572 20154
rect 13596 20102 13606 20154
rect 13606 20102 13652 20154
rect 13356 20100 13412 20102
rect 13436 20100 13492 20102
rect 13516 20100 13572 20102
rect 13596 20100 13652 20102
rect 14856 23962 14912 23964
rect 14936 23962 14992 23964
rect 15016 23962 15072 23964
rect 15096 23962 15152 23964
rect 14856 23910 14902 23962
rect 14902 23910 14912 23962
rect 14936 23910 14966 23962
rect 14966 23910 14978 23962
rect 14978 23910 14992 23962
rect 15016 23910 15030 23962
rect 15030 23910 15042 23962
rect 15042 23910 15072 23962
rect 15096 23910 15106 23962
rect 15106 23910 15152 23962
rect 14856 23908 14912 23910
rect 14936 23908 14992 23910
rect 15016 23908 15072 23910
rect 15096 23908 15152 23910
rect 15106 23588 15162 23624
rect 15106 23568 15108 23588
rect 15108 23568 15160 23588
rect 15160 23568 15162 23588
rect 14856 22874 14912 22876
rect 14936 22874 14992 22876
rect 15016 22874 15072 22876
rect 15096 22874 15152 22876
rect 14856 22822 14902 22874
rect 14902 22822 14912 22874
rect 14936 22822 14966 22874
rect 14966 22822 14978 22874
rect 14978 22822 14992 22874
rect 15016 22822 15030 22874
rect 15030 22822 15042 22874
rect 15042 22822 15072 22874
rect 15096 22822 15106 22874
rect 15106 22822 15152 22874
rect 14856 22820 14912 22822
rect 14936 22820 14992 22822
rect 15016 22820 15072 22822
rect 15096 22820 15152 22822
rect 14856 21786 14912 21788
rect 14936 21786 14992 21788
rect 15016 21786 15072 21788
rect 15096 21786 15152 21788
rect 14856 21734 14902 21786
rect 14902 21734 14912 21786
rect 14936 21734 14966 21786
rect 14966 21734 14978 21786
rect 14978 21734 14992 21786
rect 15016 21734 15030 21786
rect 15030 21734 15042 21786
rect 15042 21734 15072 21786
rect 15096 21734 15106 21786
rect 15106 21734 15152 21786
rect 14856 21732 14912 21734
rect 14936 21732 14992 21734
rect 15016 21732 15072 21734
rect 15096 21732 15152 21734
rect 15106 21004 15162 21040
rect 15106 20984 15108 21004
rect 15108 20984 15160 21004
rect 15160 20984 15162 21004
rect 14856 20698 14912 20700
rect 14936 20698 14992 20700
rect 15016 20698 15072 20700
rect 15096 20698 15152 20700
rect 14856 20646 14902 20698
rect 14902 20646 14912 20698
rect 14936 20646 14966 20698
rect 14966 20646 14978 20698
rect 14978 20646 14992 20698
rect 15016 20646 15030 20698
rect 15030 20646 15042 20698
rect 15042 20646 15072 20698
rect 15096 20646 15106 20698
rect 15106 20646 15152 20698
rect 14856 20644 14912 20646
rect 14936 20644 14992 20646
rect 15016 20644 15072 20646
rect 15096 20644 15152 20646
rect 13356 19066 13412 19068
rect 13436 19066 13492 19068
rect 13516 19066 13572 19068
rect 13596 19066 13652 19068
rect 13356 19014 13402 19066
rect 13402 19014 13412 19066
rect 13436 19014 13466 19066
rect 13466 19014 13478 19066
rect 13478 19014 13492 19066
rect 13516 19014 13530 19066
rect 13530 19014 13542 19066
rect 13542 19014 13572 19066
rect 13596 19014 13606 19066
rect 13606 19014 13652 19066
rect 13356 19012 13412 19014
rect 13436 19012 13492 19014
rect 13516 19012 13572 19014
rect 13596 19012 13652 19014
rect 13356 17978 13412 17980
rect 13436 17978 13492 17980
rect 13516 17978 13572 17980
rect 13596 17978 13652 17980
rect 13356 17926 13402 17978
rect 13402 17926 13412 17978
rect 13436 17926 13466 17978
rect 13466 17926 13478 17978
rect 13478 17926 13492 17978
rect 13516 17926 13530 17978
rect 13530 17926 13542 17978
rect 13542 17926 13572 17978
rect 13596 17926 13606 17978
rect 13606 17926 13652 17978
rect 13356 17924 13412 17926
rect 13436 17924 13492 17926
rect 13516 17924 13572 17926
rect 13596 17924 13652 17926
rect 13356 16890 13412 16892
rect 13436 16890 13492 16892
rect 13516 16890 13572 16892
rect 13596 16890 13652 16892
rect 13356 16838 13402 16890
rect 13402 16838 13412 16890
rect 13436 16838 13466 16890
rect 13466 16838 13478 16890
rect 13478 16838 13492 16890
rect 13516 16838 13530 16890
rect 13530 16838 13542 16890
rect 13542 16838 13572 16890
rect 13596 16838 13606 16890
rect 13606 16838 13652 16890
rect 13356 16836 13412 16838
rect 13436 16836 13492 16838
rect 13516 16836 13572 16838
rect 13596 16836 13652 16838
rect 13356 15802 13412 15804
rect 13436 15802 13492 15804
rect 13516 15802 13572 15804
rect 13596 15802 13652 15804
rect 13356 15750 13402 15802
rect 13402 15750 13412 15802
rect 13436 15750 13466 15802
rect 13466 15750 13478 15802
rect 13478 15750 13492 15802
rect 13516 15750 13530 15802
rect 13530 15750 13542 15802
rect 13542 15750 13572 15802
rect 13596 15750 13606 15802
rect 13606 15750 13652 15802
rect 13356 15748 13412 15750
rect 13436 15748 13492 15750
rect 13516 15748 13572 15750
rect 13596 15748 13652 15750
rect 14278 17584 14334 17640
rect 14856 19610 14912 19612
rect 14936 19610 14992 19612
rect 15016 19610 15072 19612
rect 15096 19610 15152 19612
rect 14856 19558 14902 19610
rect 14902 19558 14912 19610
rect 14936 19558 14966 19610
rect 14966 19558 14978 19610
rect 14978 19558 14992 19610
rect 15016 19558 15030 19610
rect 15030 19558 15042 19610
rect 15042 19558 15072 19610
rect 15096 19558 15106 19610
rect 15106 19558 15152 19610
rect 14856 19556 14912 19558
rect 14936 19556 14992 19558
rect 15016 19556 15072 19558
rect 15096 19556 15152 19558
rect 17856 25050 17912 25052
rect 17936 25050 17992 25052
rect 18016 25050 18072 25052
rect 18096 25050 18152 25052
rect 17856 24998 17902 25050
rect 17902 24998 17912 25050
rect 17936 24998 17966 25050
rect 17966 24998 17978 25050
rect 17978 24998 17992 25050
rect 18016 24998 18030 25050
rect 18030 24998 18042 25050
rect 18042 24998 18072 25050
rect 18096 24998 18106 25050
rect 18106 24998 18152 25050
rect 17856 24996 17912 24998
rect 17936 24996 17992 24998
rect 18016 24996 18072 24998
rect 18096 24996 18152 24998
rect 20856 25050 20912 25052
rect 20936 25050 20992 25052
rect 21016 25050 21072 25052
rect 21096 25050 21152 25052
rect 20856 24998 20902 25050
rect 20902 24998 20912 25050
rect 20936 24998 20966 25050
rect 20966 24998 20978 25050
rect 20978 24998 20992 25050
rect 21016 24998 21030 25050
rect 21030 24998 21042 25050
rect 21042 24998 21072 25050
rect 21096 24998 21106 25050
rect 21106 24998 21152 25050
rect 20856 24996 20912 24998
rect 20936 24996 20992 24998
rect 21016 24996 21072 24998
rect 21096 24996 21152 24998
rect 23856 25050 23912 25052
rect 23936 25050 23992 25052
rect 24016 25050 24072 25052
rect 24096 25050 24152 25052
rect 23856 24998 23902 25050
rect 23902 24998 23912 25050
rect 23936 24998 23966 25050
rect 23966 24998 23978 25050
rect 23978 24998 23992 25050
rect 24016 24998 24030 25050
rect 24030 24998 24042 25050
rect 24042 24998 24072 25050
rect 24096 24998 24106 25050
rect 24106 24998 24152 25050
rect 23856 24996 23912 24998
rect 23936 24996 23992 24998
rect 24016 24996 24072 24998
rect 24096 24996 24152 24998
rect 16356 24506 16412 24508
rect 16436 24506 16492 24508
rect 16516 24506 16572 24508
rect 16596 24506 16652 24508
rect 16356 24454 16402 24506
rect 16402 24454 16412 24506
rect 16436 24454 16466 24506
rect 16466 24454 16478 24506
rect 16478 24454 16492 24506
rect 16516 24454 16530 24506
rect 16530 24454 16542 24506
rect 16542 24454 16572 24506
rect 16596 24454 16606 24506
rect 16606 24454 16652 24506
rect 16356 24452 16412 24454
rect 16436 24452 16492 24454
rect 16516 24452 16572 24454
rect 16596 24452 16652 24454
rect 16356 23418 16412 23420
rect 16436 23418 16492 23420
rect 16516 23418 16572 23420
rect 16596 23418 16652 23420
rect 16356 23366 16402 23418
rect 16402 23366 16412 23418
rect 16436 23366 16466 23418
rect 16466 23366 16478 23418
rect 16478 23366 16492 23418
rect 16516 23366 16530 23418
rect 16530 23366 16542 23418
rect 16542 23366 16572 23418
rect 16596 23366 16606 23418
rect 16606 23366 16652 23418
rect 16356 23364 16412 23366
rect 16436 23364 16492 23366
rect 16516 23364 16572 23366
rect 16596 23364 16652 23366
rect 17856 23962 17912 23964
rect 17936 23962 17992 23964
rect 18016 23962 18072 23964
rect 18096 23962 18152 23964
rect 17856 23910 17902 23962
rect 17902 23910 17912 23962
rect 17936 23910 17966 23962
rect 17966 23910 17978 23962
rect 17978 23910 17992 23962
rect 18016 23910 18030 23962
rect 18030 23910 18042 23962
rect 18042 23910 18072 23962
rect 18096 23910 18106 23962
rect 18106 23910 18152 23962
rect 17856 23908 17912 23910
rect 17936 23908 17992 23910
rect 18016 23908 18072 23910
rect 18096 23908 18152 23910
rect 16356 22330 16412 22332
rect 16436 22330 16492 22332
rect 16516 22330 16572 22332
rect 16596 22330 16652 22332
rect 16356 22278 16402 22330
rect 16402 22278 16412 22330
rect 16436 22278 16466 22330
rect 16466 22278 16478 22330
rect 16478 22278 16492 22330
rect 16516 22278 16530 22330
rect 16530 22278 16542 22330
rect 16542 22278 16572 22330
rect 16596 22278 16606 22330
rect 16606 22278 16652 22330
rect 16356 22276 16412 22278
rect 16436 22276 16492 22278
rect 16516 22276 16572 22278
rect 16596 22276 16652 22278
rect 18786 23568 18842 23624
rect 17856 22874 17912 22876
rect 17936 22874 17992 22876
rect 18016 22874 18072 22876
rect 18096 22874 18152 22876
rect 17856 22822 17902 22874
rect 17902 22822 17912 22874
rect 17936 22822 17966 22874
rect 17966 22822 17978 22874
rect 17978 22822 17992 22874
rect 18016 22822 18030 22874
rect 18030 22822 18042 22874
rect 18042 22822 18072 22874
rect 18096 22822 18106 22874
rect 18106 22822 18152 22874
rect 17856 22820 17912 22822
rect 17936 22820 17992 22822
rect 18016 22820 18072 22822
rect 18096 22820 18152 22822
rect 17856 21786 17912 21788
rect 17936 21786 17992 21788
rect 18016 21786 18072 21788
rect 18096 21786 18152 21788
rect 17856 21734 17902 21786
rect 17902 21734 17912 21786
rect 17936 21734 17966 21786
rect 17966 21734 17978 21786
rect 17978 21734 17992 21786
rect 18016 21734 18030 21786
rect 18030 21734 18042 21786
rect 18042 21734 18072 21786
rect 18096 21734 18106 21786
rect 18106 21734 18152 21786
rect 17856 21732 17912 21734
rect 17936 21732 17992 21734
rect 18016 21732 18072 21734
rect 18096 21732 18152 21734
rect 14856 18522 14912 18524
rect 14936 18522 14992 18524
rect 15016 18522 15072 18524
rect 15096 18522 15152 18524
rect 14856 18470 14902 18522
rect 14902 18470 14912 18522
rect 14936 18470 14966 18522
rect 14966 18470 14978 18522
rect 14978 18470 14992 18522
rect 15016 18470 15030 18522
rect 15030 18470 15042 18522
rect 15042 18470 15072 18522
rect 15096 18470 15106 18522
rect 15106 18470 15152 18522
rect 14856 18468 14912 18470
rect 14936 18468 14992 18470
rect 15016 18468 15072 18470
rect 15096 18468 15152 18470
rect 14554 17584 14610 17640
rect 13356 14714 13412 14716
rect 13436 14714 13492 14716
rect 13516 14714 13572 14716
rect 13596 14714 13652 14716
rect 13356 14662 13402 14714
rect 13402 14662 13412 14714
rect 13436 14662 13466 14714
rect 13466 14662 13478 14714
rect 13478 14662 13492 14714
rect 13516 14662 13530 14714
rect 13530 14662 13542 14714
rect 13542 14662 13572 14714
rect 13596 14662 13606 14714
rect 13606 14662 13652 14714
rect 13356 14660 13412 14662
rect 13436 14660 13492 14662
rect 13516 14660 13572 14662
rect 13596 14660 13652 14662
rect 13726 13912 13782 13968
rect 13356 13626 13412 13628
rect 13436 13626 13492 13628
rect 13516 13626 13572 13628
rect 13596 13626 13652 13628
rect 13356 13574 13402 13626
rect 13402 13574 13412 13626
rect 13436 13574 13466 13626
rect 13466 13574 13478 13626
rect 13478 13574 13492 13626
rect 13516 13574 13530 13626
rect 13530 13574 13542 13626
rect 13542 13574 13572 13626
rect 13596 13574 13606 13626
rect 13606 13574 13652 13626
rect 13356 13572 13412 13574
rect 13436 13572 13492 13574
rect 13516 13572 13572 13574
rect 13596 13572 13652 13574
rect 11856 11994 11912 11996
rect 11936 11994 11992 11996
rect 12016 11994 12072 11996
rect 12096 11994 12152 11996
rect 11856 11942 11902 11994
rect 11902 11942 11912 11994
rect 11936 11942 11966 11994
rect 11966 11942 11978 11994
rect 11978 11942 11992 11994
rect 12016 11942 12030 11994
rect 12030 11942 12042 11994
rect 12042 11942 12072 11994
rect 12096 11942 12106 11994
rect 12106 11942 12152 11994
rect 11856 11940 11912 11942
rect 11936 11940 11992 11942
rect 12016 11940 12072 11942
rect 12096 11940 12152 11942
rect 11856 10906 11912 10908
rect 11936 10906 11992 10908
rect 12016 10906 12072 10908
rect 12096 10906 12152 10908
rect 11856 10854 11902 10906
rect 11902 10854 11912 10906
rect 11936 10854 11966 10906
rect 11966 10854 11978 10906
rect 11978 10854 11992 10906
rect 12016 10854 12030 10906
rect 12030 10854 12042 10906
rect 12042 10854 12072 10906
rect 12096 10854 12106 10906
rect 12106 10854 12152 10906
rect 11856 10852 11912 10854
rect 11936 10852 11992 10854
rect 12016 10852 12072 10854
rect 12096 10852 12152 10854
rect 11856 9818 11912 9820
rect 11936 9818 11992 9820
rect 12016 9818 12072 9820
rect 12096 9818 12152 9820
rect 11856 9766 11902 9818
rect 11902 9766 11912 9818
rect 11936 9766 11966 9818
rect 11966 9766 11978 9818
rect 11978 9766 11992 9818
rect 12016 9766 12030 9818
rect 12030 9766 12042 9818
rect 12042 9766 12072 9818
rect 12096 9766 12106 9818
rect 12106 9766 12152 9818
rect 11856 9764 11912 9766
rect 11936 9764 11992 9766
rect 12016 9764 12072 9766
rect 12096 9764 12152 9766
rect 11856 8730 11912 8732
rect 11936 8730 11992 8732
rect 12016 8730 12072 8732
rect 12096 8730 12152 8732
rect 11856 8678 11902 8730
rect 11902 8678 11912 8730
rect 11936 8678 11966 8730
rect 11966 8678 11978 8730
rect 11978 8678 11992 8730
rect 12016 8678 12030 8730
rect 12030 8678 12042 8730
rect 12042 8678 12072 8730
rect 12096 8678 12106 8730
rect 12106 8678 12152 8730
rect 11856 8676 11912 8678
rect 11936 8676 11992 8678
rect 12016 8676 12072 8678
rect 12096 8676 12152 8678
rect 11856 7642 11912 7644
rect 11936 7642 11992 7644
rect 12016 7642 12072 7644
rect 12096 7642 12152 7644
rect 11856 7590 11902 7642
rect 11902 7590 11912 7642
rect 11936 7590 11966 7642
rect 11966 7590 11978 7642
rect 11978 7590 11992 7642
rect 12016 7590 12030 7642
rect 12030 7590 12042 7642
rect 12042 7590 12072 7642
rect 12096 7590 12106 7642
rect 12106 7590 12152 7642
rect 11856 7588 11912 7590
rect 11936 7588 11992 7590
rect 12016 7588 12072 7590
rect 12096 7588 12152 7590
rect 8856 5466 8912 5468
rect 8936 5466 8992 5468
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 8856 5414 8902 5466
rect 8902 5414 8912 5466
rect 8936 5414 8966 5466
rect 8966 5414 8978 5466
rect 8978 5414 8992 5466
rect 9016 5414 9030 5466
rect 9030 5414 9042 5466
rect 9042 5414 9072 5466
rect 9096 5414 9106 5466
rect 9106 5414 9152 5466
rect 8856 5412 8912 5414
rect 8936 5412 8992 5414
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 8856 4378 8912 4380
rect 8936 4378 8992 4380
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 8856 4326 8902 4378
rect 8902 4326 8912 4378
rect 8936 4326 8966 4378
rect 8966 4326 8978 4378
rect 8978 4326 8992 4378
rect 9016 4326 9030 4378
rect 9030 4326 9042 4378
rect 9042 4326 9072 4378
rect 9096 4326 9106 4378
rect 9106 4326 9152 4378
rect 8856 4324 8912 4326
rect 8936 4324 8992 4326
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 8856 3290 8912 3292
rect 8936 3290 8992 3292
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 8856 3238 8902 3290
rect 8902 3238 8912 3290
rect 8936 3238 8966 3290
rect 8966 3238 8978 3290
rect 8978 3238 8992 3290
rect 9016 3238 9030 3290
rect 9030 3238 9042 3290
rect 9042 3238 9072 3290
rect 9096 3238 9106 3290
rect 9106 3238 9152 3290
rect 8856 3236 8912 3238
rect 8936 3236 8992 3238
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 10356 6010 10412 6012
rect 10436 6010 10492 6012
rect 10516 6010 10572 6012
rect 10596 6010 10652 6012
rect 10356 5958 10402 6010
rect 10402 5958 10412 6010
rect 10436 5958 10466 6010
rect 10466 5958 10478 6010
rect 10478 5958 10492 6010
rect 10516 5958 10530 6010
rect 10530 5958 10542 6010
rect 10542 5958 10572 6010
rect 10596 5958 10606 6010
rect 10606 5958 10652 6010
rect 10356 5956 10412 5958
rect 10436 5956 10492 5958
rect 10516 5956 10572 5958
rect 10596 5956 10652 5958
rect 10356 4922 10412 4924
rect 10436 4922 10492 4924
rect 10516 4922 10572 4924
rect 10596 4922 10652 4924
rect 10356 4870 10402 4922
rect 10402 4870 10412 4922
rect 10436 4870 10466 4922
rect 10466 4870 10478 4922
rect 10478 4870 10492 4922
rect 10516 4870 10530 4922
rect 10530 4870 10542 4922
rect 10542 4870 10572 4922
rect 10596 4870 10606 4922
rect 10606 4870 10652 4922
rect 10356 4868 10412 4870
rect 10436 4868 10492 4870
rect 10516 4868 10572 4870
rect 10596 4868 10652 4870
rect 10356 3834 10412 3836
rect 10436 3834 10492 3836
rect 10516 3834 10572 3836
rect 10596 3834 10652 3836
rect 10356 3782 10402 3834
rect 10402 3782 10412 3834
rect 10436 3782 10466 3834
rect 10466 3782 10478 3834
rect 10478 3782 10492 3834
rect 10516 3782 10530 3834
rect 10530 3782 10542 3834
rect 10542 3782 10572 3834
rect 10596 3782 10606 3834
rect 10606 3782 10652 3834
rect 10356 3780 10412 3782
rect 10436 3780 10492 3782
rect 10516 3780 10572 3782
rect 10596 3780 10652 3782
rect 11856 6554 11912 6556
rect 11936 6554 11992 6556
rect 12016 6554 12072 6556
rect 12096 6554 12152 6556
rect 11856 6502 11902 6554
rect 11902 6502 11912 6554
rect 11936 6502 11966 6554
rect 11966 6502 11978 6554
rect 11978 6502 11992 6554
rect 12016 6502 12030 6554
rect 12030 6502 12042 6554
rect 12042 6502 12072 6554
rect 12096 6502 12106 6554
rect 12106 6502 12152 6554
rect 11856 6500 11912 6502
rect 11936 6500 11992 6502
rect 12016 6500 12072 6502
rect 12096 6500 12152 6502
rect 11856 5466 11912 5468
rect 11936 5466 11992 5468
rect 12016 5466 12072 5468
rect 12096 5466 12152 5468
rect 11856 5414 11902 5466
rect 11902 5414 11912 5466
rect 11936 5414 11966 5466
rect 11966 5414 11978 5466
rect 11978 5414 11992 5466
rect 12016 5414 12030 5466
rect 12030 5414 12042 5466
rect 12042 5414 12072 5466
rect 12096 5414 12106 5466
rect 12106 5414 12152 5466
rect 11856 5412 11912 5414
rect 11936 5412 11992 5414
rect 12016 5412 12072 5414
rect 12096 5412 12152 5414
rect 11856 4378 11912 4380
rect 11936 4378 11992 4380
rect 12016 4378 12072 4380
rect 12096 4378 12152 4380
rect 11856 4326 11902 4378
rect 11902 4326 11912 4378
rect 11936 4326 11966 4378
rect 11966 4326 11978 4378
rect 11978 4326 11992 4378
rect 12016 4326 12030 4378
rect 12030 4326 12042 4378
rect 12042 4326 12072 4378
rect 12096 4326 12106 4378
rect 12106 4326 12152 4378
rect 11856 4324 11912 4326
rect 11936 4324 11992 4326
rect 12016 4324 12072 4326
rect 12096 4324 12152 4326
rect 10356 2746 10412 2748
rect 10436 2746 10492 2748
rect 10516 2746 10572 2748
rect 10596 2746 10652 2748
rect 10356 2694 10402 2746
rect 10402 2694 10412 2746
rect 10436 2694 10466 2746
rect 10466 2694 10478 2746
rect 10478 2694 10492 2746
rect 10516 2694 10530 2746
rect 10530 2694 10542 2746
rect 10542 2694 10572 2746
rect 10596 2694 10606 2746
rect 10606 2694 10652 2746
rect 10356 2692 10412 2694
rect 10436 2692 10492 2694
rect 10516 2692 10572 2694
rect 10596 2692 10652 2694
rect 11856 3290 11912 3292
rect 11936 3290 11992 3292
rect 12016 3290 12072 3292
rect 12096 3290 12152 3292
rect 11856 3238 11902 3290
rect 11902 3238 11912 3290
rect 11936 3238 11966 3290
rect 11966 3238 11978 3290
rect 11978 3238 11992 3290
rect 12016 3238 12030 3290
rect 12030 3238 12042 3290
rect 12042 3238 12072 3290
rect 12096 3238 12106 3290
rect 12106 3238 12152 3290
rect 11856 3236 11912 3238
rect 11936 3236 11992 3238
rect 12016 3236 12072 3238
rect 12096 3236 12152 3238
rect 13356 12538 13412 12540
rect 13436 12538 13492 12540
rect 13516 12538 13572 12540
rect 13596 12538 13652 12540
rect 13356 12486 13402 12538
rect 13402 12486 13412 12538
rect 13436 12486 13466 12538
rect 13466 12486 13478 12538
rect 13478 12486 13492 12538
rect 13516 12486 13530 12538
rect 13530 12486 13542 12538
rect 13542 12486 13572 12538
rect 13596 12486 13606 12538
rect 13606 12486 13652 12538
rect 13356 12484 13412 12486
rect 13436 12484 13492 12486
rect 13516 12484 13572 12486
rect 13596 12484 13652 12486
rect 14922 17584 14978 17640
rect 14856 17434 14912 17436
rect 14936 17434 14992 17436
rect 15016 17434 15072 17436
rect 15096 17434 15152 17436
rect 14856 17382 14902 17434
rect 14902 17382 14912 17434
rect 14936 17382 14966 17434
rect 14966 17382 14978 17434
rect 14978 17382 14992 17434
rect 15016 17382 15030 17434
rect 15030 17382 15042 17434
rect 15042 17382 15072 17434
rect 15096 17382 15106 17434
rect 15106 17382 15152 17434
rect 14856 17380 14912 17382
rect 14936 17380 14992 17382
rect 15016 17380 15072 17382
rect 15096 17380 15152 17382
rect 14856 16346 14912 16348
rect 14936 16346 14992 16348
rect 15016 16346 15072 16348
rect 15096 16346 15152 16348
rect 14856 16294 14902 16346
rect 14902 16294 14912 16346
rect 14936 16294 14966 16346
rect 14966 16294 14978 16346
rect 14978 16294 14992 16346
rect 15016 16294 15030 16346
rect 15030 16294 15042 16346
rect 15042 16294 15072 16346
rect 15096 16294 15106 16346
rect 15106 16294 15152 16346
rect 14856 16292 14912 16294
rect 14936 16292 14992 16294
rect 15016 16292 15072 16294
rect 15096 16292 15152 16294
rect 14856 15258 14912 15260
rect 14936 15258 14992 15260
rect 15016 15258 15072 15260
rect 15096 15258 15152 15260
rect 14856 15206 14902 15258
rect 14902 15206 14912 15258
rect 14936 15206 14966 15258
rect 14966 15206 14978 15258
rect 14978 15206 14992 15258
rect 15016 15206 15030 15258
rect 15030 15206 15042 15258
rect 15042 15206 15072 15258
rect 15096 15206 15106 15258
rect 15106 15206 15152 15258
rect 14856 15204 14912 15206
rect 14936 15204 14992 15206
rect 15016 15204 15072 15206
rect 15096 15204 15152 15206
rect 14856 14170 14912 14172
rect 14936 14170 14992 14172
rect 15016 14170 15072 14172
rect 15096 14170 15152 14172
rect 14856 14118 14902 14170
rect 14902 14118 14912 14170
rect 14936 14118 14966 14170
rect 14966 14118 14978 14170
rect 14978 14118 14992 14170
rect 15016 14118 15030 14170
rect 15030 14118 15042 14170
rect 15042 14118 15072 14170
rect 15096 14118 15106 14170
rect 15106 14118 15152 14170
rect 14856 14116 14912 14118
rect 14936 14116 14992 14118
rect 15016 14116 15072 14118
rect 15096 14116 15152 14118
rect 14856 13082 14912 13084
rect 14936 13082 14992 13084
rect 15016 13082 15072 13084
rect 15096 13082 15152 13084
rect 14856 13030 14902 13082
rect 14902 13030 14912 13082
rect 14936 13030 14966 13082
rect 14966 13030 14978 13082
rect 14978 13030 14992 13082
rect 15016 13030 15030 13082
rect 15030 13030 15042 13082
rect 15042 13030 15072 13082
rect 15096 13030 15106 13082
rect 15106 13030 15152 13082
rect 14856 13028 14912 13030
rect 14936 13028 14992 13030
rect 15016 13028 15072 13030
rect 15096 13028 15152 13030
rect 14856 11994 14912 11996
rect 14936 11994 14992 11996
rect 15016 11994 15072 11996
rect 15096 11994 15152 11996
rect 14856 11942 14902 11994
rect 14902 11942 14912 11994
rect 14936 11942 14966 11994
rect 14966 11942 14978 11994
rect 14978 11942 14992 11994
rect 15016 11942 15030 11994
rect 15030 11942 15042 11994
rect 15042 11942 15072 11994
rect 15096 11942 15106 11994
rect 15106 11942 15152 11994
rect 14856 11940 14912 11942
rect 14936 11940 14992 11942
rect 15016 11940 15072 11942
rect 15096 11940 15152 11942
rect 13356 11450 13412 11452
rect 13436 11450 13492 11452
rect 13516 11450 13572 11452
rect 13596 11450 13652 11452
rect 13356 11398 13402 11450
rect 13402 11398 13412 11450
rect 13436 11398 13466 11450
rect 13466 11398 13478 11450
rect 13478 11398 13492 11450
rect 13516 11398 13530 11450
rect 13530 11398 13542 11450
rect 13542 11398 13572 11450
rect 13596 11398 13606 11450
rect 13606 11398 13652 11450
rect 13356 11396 13412 11398
rect 13436 11396 13492 11398
rect 13516 11396 13572 11398
rect 13596 11396 13652 11398
rect 13356 10362 13412 10364
rect 13436 10362 13492 10364
rect 13516 10362 13572 10364
rect 13596 10362 13652 10364
rect 13356 10310 13402 10362
rect 13402 10310 13412 10362
rect 13436 10310 13466 10362
rect 13466 10310 13478 10362
rect 13478 10310 13492 10362
rect 13516 10310 13530 10362
rect 13530 10310 13542 10362
rect 13542 10310 13572 10362
rect 13596 10310 13606 10362
rect 13606 10310 13652 10362
rect 13356 10308 13412 10310
rect 13436 10308 13492 10310
rect 13516 10308 13572 10310
rect 13596 10308 13652 10310
rect 13356 9274 13412 9276
rect 13436 9274 13492 9276
rect 13516 9274 13572 9276
rect 13596 9274 13652 9276
rect 13356 9222 13402 9274
rect 13402 9222 13412 9274
rect 13436 9222 13466 9274
rect 13466 9222 13478 9274
rect 13478 9222 13492 9274
rect 13516 9222 13530 9274
rect 13530 9222 13542 9274
rect 13542 9222 13572 9274
rect 13596 9222 13606 9274
rect 13606 9222 13652 9274
rect 13356 9220 13412 9222
rect 13436 9220 13492 9222
rect 13516 9220 13572 9222
rect 13596 9220 13652 9222
rect 13356 8186 13412 8188
rect 13436 8186 13492 8188
rect 13516 8186 13572 8188
rect 13596 8186 13652 8188
rect 13356 8134 13402 8186
rect 13402 8134 13412 8186
rect 13436 8134 13466 8186
rect 13466 8134 13478 8186
rect 13478 8134 13492 8186
rect 13516 8134 13530 8186
rect 13530 8134 13542 8186
rect 13542 8134 13572 8186
rect 13596 8134 13606 8186
rect 13606 8134 13652 8186
rect 13356 8132 13412 8134
rect 13436 8132 13492 8134
rect 13516 8132 13572 8134
rect 13596 8132 13652 8134
rect 14370 11056 14426 11112
rect 13356 7098 13412 7100
rect 13436 7098 13492 7100
rect 13516 7098 13572 7100
rect 13596 7098 13652 7100
rect 13356 7046 13402 7098
rect 13402 7046 13412 7098
rect 13436 7046 13466 7098
rect 13466 7046 13478 7098
rect 13478 7046 13492 7098
rect 13516 7046 13530 7098
rect 13530 7046 13542 7098
rect 13542 7046 13572 7098
rect 13596 7046 13606 7098
rect 13606 7046 13652 7098
rect 13356 7044 13412 7046
rect 13436 7044 13492 7046
rect 13516 7044 13572 7046
rect 13596 7044 13652 7046
rect 13356 6010 13412 6012
rect 13436 6010 13492 6012
rect 13516 6010 13572 6012
rect 13596 6010 13652 6012
rect 13356 5958 13402 6010
rect 13402 5958 13412 6010
rect 13436 5958 13466 6010
rect 13466 5958 13478 6010
rect 13478 5958 13492 6010
rect 13516 5958 13530 6010
rect 13530 5958 13542 6010
rect 13542 5958 13572 6010
rect 13596 5958 13606 6010
rect 13606 5958 13652 6010
rect 13356 5956 13412 5958
rect 13436 5956 13492 5958
rect 13516 5956 13572 5958
rect 13596 5956 13652 5958
rect 13356 4922 13412 4924
rect 13436 4922 13492 4924
rect 13516 4922 13572 4924
rect 13596 4922 13652 4924
rect 13356 4870 13402 4922
rect 13402 4870 13412 4922
rect 13436 4870 13466 4922
rect 13466 4870 13478 4922
rect 13478 4870 13492 4922
rect 13516 4870 13530 4922
rect 13530 4870 13542 4922
rect 13542 4870 13572 4922
rect 13596 4870 13606 4922
rect 13606 4870 13652 4922
rect 13356 4868 13412 4870
rect 13436 4868 13492 4870
rect 13516 4868 13572 4870
rect 13596 4868 13652 4870
rect 13356 3834 13412 3836
rect 13436 3834 13492 3836
rect 13516 3834 13572 3836
rect 13596 3834 13652 3836
rect 13356 3782 13402 3834
rect 13402 3782 13412 3834
rect 13436 3782 13466 3834
rect 13466 3782 13478 3834
rect 13478 3782 13492 3834
rect 13516 3782 13530 3834
rect 13530 3782 13542 3834
rect 13542 3782 13572 3834
rect 13596 3782 13606 3834
rect 13606 3782 13652 3834
rect 13356 3780 13412 3782
rect 13436 3780 13492 3782
rect 13516 3780 13572 3782
rect 13596 3780 13652 3782
rect 14856 10906 14912 10908
rect 14936 10906 14992 10908
rect 15016 10906 15072 10908
rect 15096 10906 15152 10908
rect 14856 10854 14902 10906
rect 14902 10854 14912 10906
rect 14936 10854 14966 10906
rect 14966 10854 14978 10906
rect 14978 10854 14992 10906
rect 15016 10854 15030 10906
rect 15030 10854 15042 10906
rect 15042 10854 15072 10906
rect 15096 10854 15106 10906
rect 15106 10854 15152 10906
rect 14856 10852 14912 10854
rect 14936 10852 14992 10854
rect 15016 10852 15072 10854
rect 15096 10852 15152 10854
rect 14370 8336 14426 8392
rect 16356 21242 16412 21244
rect 16436 21242 16492 21244
rect 16516 21242 16572 21244
rect 16596 21242 16652 21244
rect 16356 21190 16402 21242
rect 16402 21190 16412 21242
rect 16436 21190 16466 21242
rect 16466 21190 16478 21242
rect 16478 21190 16492 21242
rect 16516 21190 16530 21242
rect 16530 21190 16542 21242
rect 16542 21190 16572 21242
rect 16596 21190 16606 21242
rect 16606 21190 16652 21242
rect 16356 21188 16412 21190
rect 16436 21188 16492 21190
rect 16516 21188 16572 21190
rect 16596 21188 16652 21190
rect 16356 20154 16412 20156
rect 16436 20154 16492 20156
rect 16516 20154 16572 20156
rect 16596 20154 16652 20156
rect 16356 20102 16402 20154
rect 16402 20102 16412 20154
rect 16436 20102 16466 20154
rect 16466 20102 16478 20154
rect 16478 20102 16492 20154
rect 16516 20102 16530 20154
rect 16530 20102 16542 20154
rect 16542 20102 16572 20154
rect 16596 20102 16606 20154
rect 16606 20102 16652 20154
rect 16356 20100 16412 20102
rect 16436 20100 16492 20102
rect 16516 20100 16572 20102
rect 16596 20100 16652 20102
rect 16356 19066 16412 19068
rect 16436 19066 16492 19068
rect 16516 19066 16572 19068
rect 16596 19066 16652 19068
rect 16356 19014 16402 19066
rect 16402 19014 16412 19066
rect 16436 19014 16466 19066
rect 16466 19014 16478 19066
rect 16478 19014 16492 19066
rect 16516 19014 16530 19066
rect 16530 19014 16542 19066
rect 16542 19014 16572 19066
rect 16596 19014 16606 19066
rect 16606 19014 16652 19066
rect 16356 19012 16412 19014
rect 16436 19012 16492 19014
rect 16516 19012 16572 19014
rect 16596 19012 16652 19014
rect 16670 18284 16726 18320
rect 19356 24506 19412 24508
rect 19436 24506 19492 24508
rect 19516 24506 19572 24508
rect 19596 24506 19652 24508
rect 19356 24454 19402 24506
rect 19402 24454 19412 24506
rect 19436 24454 19466 24506
rect 19466 24454 19478 24506
rect 19478 24454 19492 24506
rect 19516 24454 19530 24506
rect 19530 24454 19542 24506
rect 19542 24454 19572 24506
rect 19596 24454 19606 24506
rect 19606 24454 19652 24506
rect 19356 24452 19412 24454
rect 19436 24452 19492 24454
rect 19516 24452 19572 24454
rect 19596 24452 19652 24454
rect 19154 23588 19210 23624
rect 19154 23568 19156 23588
rect 19156 23568 19208 23588
rect 19208 23568 19210 23588
rect 19356 23418 19412 23420
rect 19436 23418 19492 23420
rect 19516 23418 19572 23420
rect 19596 23418 19652 23420
rect 19356 23366 19402 23418
rect 19402 23366 19412 23418
rect 19436 23366 19466 23418
rect 19466 23366 19478 23418
rect 19478 23366 19492 23418
rect 19516 23366 19530 23418
rect 19530 23366 19542 23418
rect 19542 23366 19572 23418
rect 19596 23366 19606 23418
rect 19606 23366 19652 23418
rect 19356 23364 19412 23366
rect 19436 23364 19492 23366
rect 19516 23364 19572 23366
rect 19596 23364 19652 23366
rect 19356 22330 19412 22332
rect 19436 22330 19492 22332
rect 19516 22330 19572 22332
rect 19596 22330 19652 22332
rect 19356 22278 19402 22330
rect 19402 22278 19412 22330
rect 19436 22278 19466 22330
rect 19466 22278 19478 22330
rect 19478 22278 19492 22330
rect 19516 22278 19530 22330
rect 19530 22278 19542 22330
rect 19542 22278 19572 22330
rect 19596 22278 19606 22330
rect 19606 22278 19652 22330
rect 19356 22276 19412 22278
rect 19436 22276 19492 22278
rect 19516 22276 19572 22278
rect 19596 22276 19652 22278
rect 17856 20698 17912 20700
rect 17936 20698 17992 20700
rect 18016 20698 18072 20700
rect 18096 20698 18152 20700
rect 17856 20646 17902 20698
rect 17902 20646 17912 20698
rect 17936 20646 17966 20698
rect 17966 20646 17978 20698
rect 17978 20646 17992 20698
rect 18016 20646 18030 20698
rect 18030 20646 18042 20698
rect 18042 20646 18072 20698
rect 18096 20646 18106 20698
rect 18106 20646 18152 20698
rect 17856 20644 17912 20646
rect 17936 20644 17992 20646
rect 18016 20644 18072 20646
rect 18096 20644 18152 20646
rect 16670 18264 16672 18284
rect 16672 18264 16724 18284
rect 16724 18264 16726 18284
rect 16356 17978 16412 17980
rect 16436 17978 16492 17980
rect 16516 17978 16572 17980
rect 16596 17978 16652 17980
rect 16356 17926 16402 17978
rect 16402 17926 16412 17978
rect 16436 17926 16466 17978
rect 16466 17926 16478 17978
rect 16478 17926 16492 17978
rect 16516 17926 16530 17978
rect 16530 17926 16542 17978
rect 16542 17926 16572 17978
rect 16596 17926 16606 17978
rect 16606 17926 16652 17978
rect 16356 17924 16412 17926
rect 16436 17924 16492 17926
rect 16516 17924 16572 17926
rect 16596 17924 16652 17926
rect 16356 16890 16412 16892
rect 16436 16890 16492 16892
rect 16516 16890 16572 16892
rect 16596 16890 16652 16892
rect 16356 16838 16402 16890
rect 16402 16838 16412 16890
rect 16436 16838 16466 16890
rect 16466 16838 16478 16890
rect 16478 16838 16492 16890
rect 16516 16838 16530 16890
rect 16530 16838 16542 16890
rect 16542 16838 16572 16890
rect 16596 16838 16606 16890
rect 16606 16838 16652 16890
rect 16356 16836 16412 16838
rect 16436 16836 16492 16838
rect 16516 16836 16572 16838
rect 16596 16836 16652 16838
rect 16356 15802 16412 15804
rect 16436 15802 16492 15804
rect 16516 15802 16572 15804
rect 16596 15802 16652 15804
rect 16356 15750 16402 15802
rect 16402 15750 16412 15802
rect 16436 15750 16466 15802
rect 16466 15750 16478 15802
rect 16478 15750 16492 15802
rect 16516 15750 16530 15802
rect 16530 15750 16542 15802
rect 16542 15750 16572 15802
rect 16596 15750 16606 15802
rect 16606 15750 16652 15802
rect 16356 15748 16412 15750
rect 16436 15748 16492 15750
rect 16516 15748 16572 15750
rect 16596 15748 16652 15750
rect 19356 21242 19412 21244
rect 19436 21242 19492 21244
rect 19516 21242 19572 21244
rect 19596 21242 19652 21244
rect 19356 21190 19402 21242
rect 19402 21190 19412 21242
rect 19436 21190 19466 21242
rect 19466 21190 19478 21242
rect 19478 21190 19492 21242
rect 19516 21190 19530 21242
rect 19530 21190 19542 21242
rect 19542 21190 19572 21242
rect 19596 21190 19606 21242
rect 19606 21190 19652 21242
rect 19356 21188 19412 21190
rect 19436 21188 19492 21190
rect 19516 21188 19572 21190
rect 19596 21188 19652 21190
rect 19356 20154 19412 20156
rect 19436 20154 19492 20156
rect 19516 20154 19572 20156
rect 19596 20154 19652 20156
rect 19356 20102 19402 20154
rect 19402 20102 19412 20154
rect 19436 20102 19466 20154
rect 19466 20102 19478 20154
rect 19478 20102 19492 20154
rect 19516 20102 19530 20154
rect 19530 20102 19542 20154
rect 19542 20102 19572 20154
rect 19596 20102 19606 20154
rect 19606 20102 19652 20154
rect 19356 20100 19412 20102
rect 19436 20100 19492 20102
rect 19516 20100 19572 20102
rect 19596 20100 19652 20102
rect 17856 19610 17912 19612
rect 17936 19610 17992 19612
rect 18016 19610 18072 19612
rect 18096 19610 18152 19612
rect 17856 19558 17902 19610
rect 17902 19558 17912 19610
rect 17936 19558 17966 19610
rect 17966 19558 17978 19610
rect 17978 19558 17992 19610
rect 18016 19558 18030 19610
rect 18030 19558 18042 19610
rect 18042 19558 18072 19610
rect 18096 19558 18106 19610
rect 18106 19558 18152 19610
rect 17856 19556 17912 19558
rect 17936 19556 17992 19558
rect 18016 19556 18072 19558
rect 18096 19556 18152 19558
rect 17856 18522 17912 18524
rect 17936 18522 17992 18524
rect 18016 18522 18072 18524
rect 18096 18522 18152 18524
rect 17856 18470 17902 18522
rect 17902 18470 17912 18522
rect 17936 18470 17966 18522
rect 17966 18470 17978 18522
rect 17978 18470 17992 18522
rect 18016 18470 18030 18522
rect 18030 18470 18042 18522
rect 18042 18470 18072 18522
rect 18096 18470 18106 18522
rect 18106 18470 18152 18522
rect 17856 18468 17912 18470
rect 17936 18468 17992 18470
rect 18016 18468 18072 18470
rect 18096 18468 18152 18470
rect 19356 19066 19412 19068
rect 19436 19066 19492 19068
rect 19516 19066 19572 19068
rect 19596 19066 19652 19068
rect 19356 19014 19402 19066
rect 19402 19014 19412 19066
rect 19436 19014 19466 19066
rect 19466 19014 19478 19066
rect 19478 19014 19492 19066
rect 19516 19014 19530 19066
rect 19530 19014 19542 19066
rect 19542 19014 19572 19066
rect 19596 19014 19606 19066
rect 19606 19014 19652 19066
rect 19356 19012 19412 19014
rect 19436 19012 19492 19014
rect 19516 19012 19572 19014
rect 19596 19012 19652 19014
rect 17856 17434 17912 17436
rect 17936 17434 17992 17436
rect 18016 17434 18072 17436
rect 18096 17434 18152 17436
rect 17856 17382 17902 17434
rect 17902 17382 17912 17434
rect 17936 17382 17966 17434
rect 17966 17382 17978 17434
rect 17978 17382 17992 17434
rect 18016 17382 18030 17434
rect 18030 17382 18042 17434
rect 18042 17382 18072 17434
rect 18096 17382 18106 17434
rect 18106 17382 18152 17434
rect 17856 17380 17912 17382
rect 17936 17380 17992 17382
rect 18016 17380 18072 17382
rect 18096 17380 18152 17382
rect 17856 16346 17912 16348
rect 17936 16346 17992 16348
rect 18016 16346 18072 16348
rect 18096 16346 18152 16348
rect 17856 16294 17902 16346
rect 17902 16294 17912 16346
rect 17936 16294 17966 16346
rect 17966 16294 17978 16346
rect 17978 16294 17992 16346
rect 18016 16294 18030 16346
rect 18030 16294 18042 16346
rect 18042 16294 18072 16346
rect 18096 16294 18106 16346
rect 18106 16294 18152 16346
rect 17856 16292 17912 16294
rect 17936 16292 17992 16294
rect 18016 16292 18072 16294
rect 18096 16292 18152 16294
rect 16356 14714 16412 14716
rect 16436 14714 16492 14716
rect 16516 14714 16572 14716
rect 16596 14714 16652 14716
rect 16356 14662 16402 14714
rect 16402 14662 16412 14714
rect 16436 14662 16466 14714
rect 16466 14662 16478 14714
rect 16478 14662 16492 14714
rect 16516 14662 16530 14714
rect 16530 14662 16542 14714
rect 16542 14662 16572 14714
rect 16596 14662 16606 14714
rect 16606 14662 16652 14714
rect 16356 14660 16412 14662
rect 16436 14660 16492 14662
rect 16516 14660 16572 14662
rect 16596 14660 16652 14662
rect 16356 13626 16412 13628
rect 16436 13626 16492 13628
rect 16516 13626 16572 13628
rect 16596 13626 16652 13628
rect 16356 13574 16402 13626
rect 16402 13574 16412 13626
rect 16436 13574 16466 13626
rect 16466 13574 16478 13626
rect 16478 13574 16492 13626
rect 16516 13574 16530 13626
rect 16530 13574 16542 13626
rect 16542 13574 16572 13626
rect 16596 13574 16606 13626
rect 16606 13574 16652 13626
rect 16356 13572 16412 13574
rect 16436 13572 16492 13574
rect 16516 13572 16572 13574
rect 16596 13572 16652 13574
rect 14856 9818 14912 9820
rect 14936 9818 14992 9820
rect 15016 9818 15072 9820
rect 15096 9818 15152 9820
rect 14856 9766 14902 9818
rect 14902 9766 14912 9818
rect 14936 9766 14966 9818
rect 14966 9766 14978 9818
rect 14978 9766 14992 9818
rect 15016 9766 15030 9818
rect 15030 9766 15042 9818
rect 15042 9766 15072 9818
rect 15096 9766 15106 9818
rect 15106 9766 15152 9818
rect 14856 9764 14912 9766
rect 14936 9764 14992 9766
rect 15016 9764 15072 9766
rect 15096 9764 15152 9766
rect 14856 8730 14912 8732
rect 14936 8730 14992 8732
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 14856 8678 14902 8730
rect 14902 8678 14912 8730
rect 14936 8678 14966 8730
rect 14966 8678 14978 8730
rect 14978 8678 14992 8730
rect 15016 8678 15030 8730
rect 15030 8678 15042 8730
rect 15042 8678 15072 8730
rect 15096 8678 15106 8730
rect 15106 8678 15152 8730
rect 14856 8676 14912 8678
rect 14936 8676 14992 8678
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 16356 12538 16412 12540
rect 16436 12538 16492 12540
rect 16516 12538 16572 12540
rect 16596 12538 16652 12540
rect 16356 12486 16402 12538
rect 16402 12486 16412 12538
rect 16436 12486 16466 12538
rect 16466 12486 16478 12538
rect 16478 12486 16492 12538
rect 16516 12486 16530 12538
rect 16530 12486 16542 12538
rect 16542 12486 16572 12538
rect 16596 12486 16606 12538
rect 16606 12486 16652 12538
rect 16356 12484 16412 12486
rect 16436 12484 16492 12486
rect 16516 12484 16572 12486
rect 16596 12484 16652 12486
rect 16356 11450 16412 11452
rect 16436 11450 16492 11452
rect 16516 11450 16572 11452
rect 16596 11450 16652 11452
rect 16356 11398 16402 11450
rect 16402 11398 16412 11450
rect 16436 11398 16466 11450
rect 16466 11398 16478 11450
rect 16478 11398 16492 11450
rect 16516 11398 16530 11450
rect 16530 11398 16542 11450
rect 16542 11398 16572 11450
rect 16596 11398 16606 11450
rect 16606 11398 16652 11450
rect 16356 11396 16412 11398
rect 16436 11396 16492 11398
rect 16516 11396 16572 11398
rect 16596 11396 16652 11398
rect 16356 10362 16412 10364
rect 16436 10362 16492 10364
rect 16516 10362 16572 10364
rect 16596 10362 16652 10364
rect 16356 10310 16402 10362
rect 16402 10310 16412 10362
rect 16436 10310 16466 10362
rect 16466 10310 16478 10362
rect 16478 10310 16492 10362
rect 16516 10310 16530 10362
rect 16530 10310 16542 10362
rect 16542 10310 16572 10362
rect 16596 10310 16606 10362
rect 16606 10310 16652 10362
rect 16356 10308 16412 10310
rect 16436 10308 16492 10310
rect 16516 10308 16572 10310
rect 16596 10308 16652 10310
rect 16356 9274 16412 9276
rect 16436 9274 16492 9276
rect 16516 9274 16572 9276
rect 16596 9274 16652 9276
rect 16356 9222 16402 9274
rect 16402 9222 16412 9274
rect 16436 9222 16466 9274
rect 16466 9222 16478 9274
rect 16478 9222 16492 9274
rect 16516 9222 16530 9274
rect 16530 9222 16542 9274
rect 16542 9222 16572 9274
rect 16596 9222 16606 9274
rect 16606 9222 16652 9274
rect 16356 9220 16412 9222
rect 16436 9220 16492 9222
rect 16516 9220 16572 9222
rect 16596 9220 16652 9222
rect 17856 15258 17912 15260
rect 17936 15258 17992 15260
rect 18016 15258 18072 15260
rect 18096 15258 18152 15260
rect 17856 15206 17902 15258
rect 17902 15206 17912 15258
rect 17936 15206 17966 15258
rect 17966 15206 17978 15258
rect 17978 15206 17992 15258
rect 18016 15206 18030 15258
rect 18030 15206 18042 15258
rect 18042 15206 18072 15258
rect 18096 15206 18106 15258
rect 18106 15206 18152 15258
rect 17856 15204 17912 15206
rect 17936 15204 17992 15206
rect 18016 15204 18072 15206
rect 18096 15204 18152 15206
rect 22356 24506 22412 24508
rect 22436 24506 22492 24508
rect 22516 24506 22572 24508
rect 22596 24506 22652 24508
rect 22356 24454 22402 24506
rect 22402 24454 22412 24506
rect 22436 24454 22466 24506
rect 22466 24454 22478 24506
rect 22478 24454 22492 24506
rect 22516 24454 22530 24506
rect 22530 24454 22542 24506
rect 22542 24454 22572 24506
rect 22596 24454 22606 24506
rect 22606 24454 22652 24506
rect 22356 24452 22412 24454
rect 22436 24452 22492 24454
rect 22516 24452 22572 24454
rect 22596 24452 22652 24454
rect 20856 23962 20912 23964
rect 20936 23962 20992 23964
rect 21016 23962 21072 23964
rect 21096 23962 21152 23964
rect 20856 23910 20902 23962
rect 20902 23910 20912 23962
rect 20936 23910 20966 23962
rect 20966 23910 20978 23962
rect 20978 23910 20992 23962
rect 21016 23910 21030 23962
rect 21030 23910 21042 23962
rect 21042 23910 21072 23962
rect 21096 23910 21106 23962
rect 21106 23910 21152 23962
rect 20856 23908 20912 23910
rect 20936 23908 20992 23910
rect 21016 23908 21072 23910
rect 21096 23908 21152 23910
rect 23856 23962 23912 23964
rect 23936 23962 23992 23964
rect 24016 23962 24072 23964
rect 24096 23962 24152 23964
rect 23856 23910 23902 23962
rect 23902 23910 23912 23962
rect 23936 23910 23966 23962
rect 23966 23910 23978 23962
rect 23978 23910 23992 23962
rect 24016 23910 24030 23962
rect 24030 23910 24042 23962
rect 24042 23910 24072 23962
rect 24096 23910 24106 23962
rect 24106 23910 24152 23962
rect 23856 23908 23912 23910
rect 23936 23908 23992 23910
rect 24016 23908 24072 23910
rect 24096 23908 24152 23910
rect 22356 23418 22412 23420
rect 22436 23418 22492 23420
rect 22516 23418 22572 23420
rect 22596 23418 22652 23420
rect 22356 23366 22402 23418
rect 22402 23366 22412 23418
rect 22436 23366 22466 23418
rect 22466 23366 22478 23418
rect 22478 23366 22492 23418
rect 22516 23366 22530 23418
rect 22530 23366 22542 23418
rect 22542 23366 22572 23418
rect 22596 23366 22606 23418
rect 22606 23366 22652 23418
rect 22356 23364 22412 23366
rect 22436 23364 22492 23366
rect 22516 23364 22572 23366
rect 22596 23364 22652 23366
rect 20856 22874 20912 22876
rect 20936 22874 20992 22876
rect 21016 22874 21072 22876
rect 21096 22874 21152 22876
rect 20856 22822 20902 22874
rect 20902 22822 20912 22874
rect 20936 22822 20966 22874
rect 20966 22822 20978 22874
rect 20978 22822 20992 22874
rect 21016 22822 21030 22874
rect 21030 22822 21042 22874
rect 21042 22822 21072 22874
rect 21096 22822 21106 22874
rect 21106 22822 21152 22874
rect 20856 22820 20912 22822
rect 20936 22820 20992 22822
rect 21016 22820 21072 22822
rect 21096 22820 21152 22822
rect 23856 22874 23912 22876
rect 23936 22874 23992 22876
rect 24016 22874 24072 22876
rect 24096 22874 24152 22876
rect 23856 22822 23902 22874
rect 23902 22822 23912 22874
rect 23936 22822 23966 22874
rect 23966 22822 23978 22874
rect 23978 22822 23992 22874
rect 24016 22822 24030 22874
rect 24030 22822 24042 22874
rect 24042 22822 24072 22874
rect 24096 22822 24106 22874
rect 24106 22822 24152 22874
rect 23856 22820 23912 22822
rect 23936 22820 23992 22822
rect 24016 22820 24072 22822
rect 24096 22820 24152 22822
rect 22356 22330 22412 22332
rect 22436 22330 22492 22332
rect 22516 22330 22572 22332
rect 22596 22330 22652 22332
rect 22356 22278 22402 22330
rect 22402 22278 22412 22330
rect 22436 22278 22466 22330
rect 22466 22278 22478 22330
rect 22478 22278 22492 22330
rect 22516 22278 22530 22330
rect 22530 22278 22542 22330
rect 22542 22278 22572 22330
rect 22596 22278 22606 22330
rect 22606 22278 22652 22330
rect 22356 22276 22412 22278
rect 22436 22276 22492 22278
rect 22516 22276 22572 22278
rect 22596 22276 22652 22278
rect 20856 21786 20912 21788
rect 20936 21786 20992 21788
rect 21016 21786 21072 21788
rect 21096 21786 21152 21788
rect 20856 21734 20902 21786
rect 20902 21734 20912 21786
rect 20936 21734 20966 21786
rect 20966 21734 20978 21786
rect 20978 21734 20992 21786
rect 21016 21734 21030 21786
rect 21030 21734 21042 21786
rect 21042 21734 21072 21786
rect 21096 21734 21106 21786
rect 21106 21734 21152 21786
rect 20856 21732 20912 21734
rect 20936 21732 20992 21734
rect 21016 21732 21072 21734
rect 21096 21732 21152 21734
rect 23856 21786 23912 21788
rect 23936 21786 23992 21788
rect 24016 21786 24072 21788
rect 24096 21786 24152 21788
rect 23856 21734 23902 21786
rect 23902 21734 23912 21786
rect 23936 21734 23966 21786
rect 23966 21734 23978 21786
rect 23978 21734 23992 21786
rect 24016 21734 24030 21786
rect 24030 21734 24042 21786
rect 24042 21734 24072 21786
rect 24096 21734 24106 21786
rect 24106 21734 24152 21786
rect 23856 21732 23912 21734
rect 23936 21732 23992 21734
rect 24016 21732 24072 21734
rect 24096 21732 24152 21734
rect 20856 20698 20912 20700
rect 20936 20698 20992 20700
rect 21016 20698 21072 20700
rect 21096 20698 21152 20700
rect 20856 20646 20902 20698
rect 20902 20646 20912 20698
rect 20936 20646 20966 20698
rect 20966 20646 20978 20698
rect 20978 20646 20992 20698
rect 21016 20646 21030 20698
rect 21030 20646 21042 20698
rect 21042 20646 21072 20698
rect 21096 20646 21106 20698
rect 21106 20646 21152 20698
rect 20856 20644 20912 20646
rect 20936 20644 20992 20646
rect 21016 20644 21072 20646
rect 21096 20644 21152 20646
rect 22356 21242 22412 21244
rect 22436 21242 22492 21244
rect 22516 21242 22572 21244
rect 22596 21242 22652 21244
rect 22356 21190 22402 21242
rect 22402 21190 22412 21242
rect 22436 21190 22466 21242
rect 22466 21190 22478 21242
rect 22478 21190 22492 21242
rect 22516 21190 22530 21242
rect 22530 21190 22542 21242
rect 22542 21190 22572 21242
rect 22596 21190 22606 21242
rect 22606 21190 22652 21242
rect 22356 21188 22412 21190
rect 22436 21188 22492 21190
rect 22516 21188 22572 21190
rect 22596 21188 22652 21190
rect 23570 21120 23626 21176
rect 20856 19610 20912 19612
rect 20936 19610 20992 19612
rect 21016 19610 21072 19612
rect 21096 19610 21152 19612
rect 20856 19558 20902 19610
rect 20902 19558 20912 19610
rect 20936 19558 20966 19610
rect 20966 19558 20978 19610
rect 20978 19558 20992 19610
rect 21016 19558 21030 19610
rect 21030 19558 21042 19610
rect 21042 19558 21072 19610
rect 21096 19558 21106 19610
rect 21106 19558 21152 19610
rect 20856 19556 20912 19558
rect 20936 19556 20992 19558
rect 21016 19556 21072 19558
rect 21096 19556 21152 19558
rect 19356 17978 19412 17980
rect 19436 17978 19492 17980
rect 19516 17978 19572 17980
rect 19596 17978 19652 17980
rect 19356 17926 19402 17978
rect 19402 17926 19412 17978
rect 19436 17926 19466 17978
rect 19466 17926 19478 17978
rect 19478 17926 19492 17978
rect 19516 17926 19530 17978
rect 19530 17926 19542 17978
rect 19542 17926 19572 17978
rect 19596 17926 19606 17978
rect 19606 17926 19652 17978
rect 19356 17924 19412 17926
rect 19436 17924 19492 17926
rect 19516 17924 19572 17926
rect 19596 17924 19652 17926
rect 20856 18522 20912 18524
rect 20936 18522 20992 18524
rect 21016 18522 21072 18524
rect 21096 18522 21152 18524
rect 20856 18470 20902 18522
rect 20902 18470 20912 18522
rect 20936 18470 20966 18522
rect 20966 18470 20978 18522
rect 20978 18470 20992 18522
rect 21016 18470 21030 18522
rect 21030 18470 21042 18522
rect 21042 18470 21072 18522
rect 21096 18470 21106 18522
rect 21106 18470 21152 18522
rect 20856 18468 20912 18470
rect 20936 18468 20992 18470
rect 21016 18468 21072 18470
rect 21096 18468 21152 18470
rect 20718 17856 20774 17912
rect 19356 16890 19412 16892
rect 19436 16890 19492 16892
rect 19516 16890 19572 16892
rect 19596 16890 19652 16892
rect 19356 16838 19402 16890
rect 19402 16838 19412 16890
rect 19436 16838 19466 16890
rect 19466 16838 19478 16890
rect 19478 16838 19492 16890
rect 19516 16838 19530 16890
rect 19530 16838 19542 16890
rect 19542 16838 19572 16890
rect 19596 16838 19606 16890
rect 19606 16838 19652 16890
rect 19356 16836 19412 16838
rect 19436 16836 19492 16838
rect 19516 16836 19572 16838
rect 19596 16836 19652 16838
rect 20856 17434 20912 17436
rect 20936 17434 20992 17436
rect 21016 17434 21072 17436
rect 21096 17434 21152 17436
rect 20856 17382 20902 17434
rect 20902 17382 20912 17434
rect 20936 17382 20966 17434
rect 20966 17382 20978 17434
rect 20978 17382 20992 17434
rect 21016 17382 21030 17434
rect 21030 17382 21042 17434
rect 21042 17382 21072 17434
rect 21096 17382 21106 17434
rect 21106 17382 21152 17434
rect 20856 17380 20912 17382
rect 20936 17380 20992 17382
rect 21016 17380 21072 17382
rect 21096 17380 21152 17382
rect 23856 20698 23912 20700
rect 23936 20698 23992 20700
rect 24016 20698 24072 20700
rect 24096 20698 24152 20700
rect 23856 20646 23902 20698
rect 23902 20646 23912 20698
rect 23936 20646 23966 20698
rect 23966 20646 23978 20698
rect 23978 20646 23992 20698
rect 24016 20646 24030 20698
rect 24030 20646 24042 20698
rect 24042 20646 24072 20698
rect 24096 20646 24106 20698
rect 24106 20646 24152 20698
rect 23856 20644 23912 20646
rect 23936 20644 23992 20646
rect 24016 20644 24072 20646
rect 24096 20644 24152 20646
rect 20856 16346 20912 16348
rect 20936 16346 20992 16348
rect 21016 16346 21072 16348
rect 21096 16346 21152 16348
rect 20856 16294 20902 16346
rect 20902 16294 20912 16346
rect 20936 16294 20966 16346
rect 20966 16294 20978 16346
rect 20978 16294 20992 16346
rect 21016 16294 21030 16346
rect 21030 16294 21042 16346
rect 21042 16294 21072 16346
rect 21096 16294 21106 16346
rect 21106 16294 21152 16346
rect 20856 16292 20912 16294
rect 20936 16292 20992 16294
rect 21016 16292 21072 16294
rect 21096 16292 21152 16294
rect 19356 15802 19412 15804
rect 19436 15802 19492 15804
rect 19516 15802 19572 15804
rect 19596 15802 19652 15804
rect 19356 15750 19402 15802
rect 19402 15750 19412 15802
rect 19436 15750 19466 15802
rect 19466 15750 19478 15802
rect 19478 15750 19492 15802
rect 19516 15750 19530 15802
rect 19530 15750 19542 15802
rect 19542 15750 19572 15802
rect 19596 15750 19606 15802
rect 19606 15750 19652 15802
rect 19356 15748 19412 15750
rect 19436 15748 19492 15750
rect 19516 15748 19572 15750
rect 19596 15748 19652 15750
rect 19246 15580 19248 15600
rect 19248 15580 19300 15600
rect 19300 15580 19302 15600
rect 19246 15544 19302 15580
rect 17856 14170 17912 14172
rect 17936 14170 17992 14172
rect 18016 14170 18072 14172
rect 18096 14170 18152 14172
rect 17856 14118 17902 14170
rect 17902 14118 17912 14170
rect 17936 14118 17966 14170
rect 17966 14118 17978 14170
rect 17978 14118 17992 14170
rect 18016 14118 18030 14170
rect 18030 14118 18042 14170
rect 18042 14118 18072 14170
rect 18096 14118 18106 14170
rect 18106 14118 18152 14170
rect 17856 14116 17912 14118
rect 17936 14116 17992 14118
rect 18016 14116 18072 14118
rect 18096 14116 18152 14118
rect 19356 14714 19412 14716
rect 19436 14714 19492 14716
rect 19516 14714 19572 14716
rect 19596 14714 19652 14716
rect 19356 14662 19402 14714
rect 19402 14662 19412 14714
rect 19436 14662 19466 14714
rect 19466 14662 19478 14714
rect 19478 14662 19492 14714
rect 19516 14662 19530 14714
rect 19530 14662 19542 14714
rect 19542 14662 19572 14714
rect 19596 14662 19606 14714
rect 19606 14662 19652 14714
rect 19356 14660 19412 14662
rect 19436 14660 19492 14662
rect 19516 14660 19572 14662
rect 19596 14660 19652 14662
rect 17856 13082 17912 13084
rect 17936 13082 17992 13084
rect 18016 13082 18072 13084
rect 18096 13082 18152 13084
rect 17856 13030 17902 13082
rect 17902 13030 17912 13082
rect 17936 13030 17966 13082
rect 17966 13030 17978 13082
rect 17978 13030 17992 13082
rect 18016 13030 18030 13082
rect 18030 13030 18042 13082
rect 18042 13030 18072 13082
rect 18096 13030 18106 13082
rect 18106 13030 18152 13082
rect 17856 13028 17912 13030
rect 17936 13028 17992 13030
rect 18016 13028 18072 13030
rect 18096 13028 18152 13030
rect 17856 11994 17912 11996
rect 17936 11994 17992 11996
rect 18016 11994 18072 11996
rect 18096 11994 18152 11996
rect 17856 11942 17902 11994
rect 17902 11942 17912 11994
rect 17936 11942 17966 11994
rect 17966 11942 17978 11994
rect 17978 11942 17992 11994
rect 18016 11942 18030 11994
rect 18030 11942 18042 11994
rect 18042 11942 18072 11994
rect 18096 11942 18106 11994
rect 18106 11942 18152 11994
rect 17856 11940 17912 11942
rect 17936 11940 17992 11942
rect 18016 11940 18072 11942
rect 18096 11940 18152 11942
rect 19356 13626 19412 13628
rect 19436 13626 19492 13628
rect 19516 13626 19572 13628
rect 19596 13626 19652 13628
rect 19356 13574 19402 13626
rect 19402 13574 19412 13626
rect 19436 13574 19466 13626
rect 19466 13574 19478 13626
rect 19478 13574 19492 13626
rect 19516 13574 19530 13626
rect 19530 13574 19542 13626
rect 19542 13574 19572 13626
rect 19596 13574 19606 13626
rect 19606 13574 19652 13626
rect 19356 13572 19412 13574
rect 19436 13572 19492 13574
rect 19516 13572 19572 13574
rect 19596 13572 19652 13574
rect 20856 15258 20912 15260
rect 20936 15258 20992 15260
rect 21016 15258 21072 15260
rect 21096 15258 21152 15260
rect 20856 15206 20902 15258
rect 20902 15206 20912 15258
rect 20936 15206 20966 15258
rect 20966 15206 20978 15258
rect 20978 15206 20992 15258
rect 21016 15206 21030 15258
rect 21030 15206 21042 15258
rect 21042 15206 21072 15258
rect 21096 15206 21106 15258
rect 21106 15206 21152 15258
rect 20856 15204 20912 15206
rect 20936 15204 20992 15206
rect 21016 15204 21072 15206
rect 21096 15204 21152 15206
rect 21546 15000 21602 15056
rect 20856 14170 20912 14172
rect 20936 14170 20992 14172
rect 21016 14170 21072 14172
rect 21096 14170 21152 14172
rect 20856 14118 20902 14170
rect 20902 14118 20912 14170
rect 20936 14118 20966 14170
rect 20966 14118 20978 14170
rect 20978 14118 20992 14170
rect 21016 14118 21030 14170
rect 21030 14118 21042 14170
rect 21042 14118 21072 14170
rect 21096 14118 21106 14170
rect 21106 14118 21152 14170
rect 20856 14116 20912 14118
rect 20936 14116 20992 14118
rect 21016 14116 21072 14118
rect 21096 14116 21152 14118
rect 19356 12538 19412 12540
rect 19436 12538 19492 12540
rect 19516 12538 19572 12540
rect 19596 12538 19652 12540
rect 19356 12486 19402 12538
rect 19402 12486 19412 12538
rect 19436 12486 19466 12538
rect 19466 12486 19478 12538
rect 19478 12486 19492 12538
rect 19516 12486 19530 12538
rect 19530 12486 19542 12538
rect 19542 12486 19572 12538
rect 19596 12486 19606 12538
rect 19606 12486 19652 12538
rect 19356 12484 19412 12486
rect 19436 12484 19492 12486
rect 19516 12484 19572 12486
rect 19596 12484 19652 12486
rect 19356 11450 19412 11452
rect 19436 11450 19492 11452
rect 19516 11450 19572 11452
rect 19596 11450 19652 11452
rect 19356 11398 19402 11450
rect 19402 11398 19412 11450
rect 19436 11398 19466 11450
rect 19466 11398 19478 11450
rect 19478 11398 19492 11450
rect 19516 11398 19530 11450
rect 19530 11398 19542 11450
rect 19542 11398 19572 11450
rect 19596 11398 19606 11450
rect 19606 11398 19652 11450
rect 19356 11396 19412 11398
rect 19436 11396 19492 11398
rect 19516 11396 19572 11398
rect 19596 11396 19652 11398
rect 20856 13082 20912 13084
rect 20936 13082 20992 13084
rect 21016 13082 21072 13084
rect 21096 13082 21152 13084
rect 20856 13030 20902 13082
rect 20902 13030 20912 13082
rect 20936 13030 20966 13082
rect 20966 13030 20978 13082
rect 20978 13030 20992 13082
rect 21016 13030 21030 13082
rect 21030 13030 21042 13082
rect 21042 13030 21072 13082
rect 21096 13030 21106 13082
rect 21106 13030 21152 13082
rect 20856 13028 20912 13030
rect 20936 13028 20992 13030
rect 21016 13028 21072 13030
rect 21096 13028 21152 13030
rect 22356 20154 22412 20156
rect 22436 20154 22492 20156
rect 22516 20154 22572 20156
rect 22596 20154 22652 20156
rect 22356 20102 22402 20154
rect 22402 20102 22412 20154
rect 22436 20102 22466 20154
rect 22466 20102 22478 20154
rect 22478 20102 22492 20154
rect 22516 20102 22530 20154
rect 22530 20102 22542 20154
rect 22542 20102 22572 20154
rect 22596 20102 22606 20154
rect 22606 20102 22652 20154
rect 22356 20100 22412 20102
rect 22436 20100 22492 20102
rect 22516 20100 22572 20102
rect 22596 20100 22652 20102
rect 22356 19066 22412 19068
rect 22436 19066 22492 19068
rect 22516 19066 22572 19068
rect 22596 19066 22652 19068
rect 22356 19014 22402 19066
rect 22402 19014 22412 19066
rect 22436 19014 22466 19066
rect 22466 19014 22478 19066
rect 22478 19014 22492 19066
rect 22516 19014 22530 19066
rect 22530 19014 22542 19066
rect 22542 19014 22572 19066
rect 22596 19014 22606 19066
rect 22606 19014 22652 19066
rect 22356 19012 22412 19014
rect 22436 19012 22492 19014
rect 22516 19012 22572 19014
rect 22596 19012 22652 19014
rect 22374 18128 22430 18184
rect 22356 17978 22412 17980
rect 22436 17978 22492 17980
rect 22516 17978 22572 17980
rect 22596 17978 22652 17980
rect 22356 17926 22402 17978
rect 22402 17926 22412 17978
rect 22436 17926 22466 17978
rect 22466 17926 22478 17978
rect 22478 17926 22492 17978
rect 22516 17926 22530 17978
rect 22530 17926 22542 17978
rect 22542 17926 22572 17978
rect 22596 17926 22606 17978
rect 22606 17926 22652 17978
rect 22356 17924 22412 17926
rect 22436 17924 22492 17926
rect 22516 17924 22572 17926
rect 22596 17924 22652 17926
rect 22356 16890 22412 16892
rect 22436 16890 22492 16892
rect 22516 16890 22572 16892
rect 22596 16890 22652 16892
rect 22356 16838 22402 16890
rect 22402 16838 22412 16890
rect 22436 16838 22466 16890
rect 22466 16838 22478 16890
rect 22478 16838 22492 16890
rect 22516 16838 22530 16890
rect 22530 16838 22542 16890
rect 22542 16838 22572 16890
rect 22596 16838 22606 16890
rect 22606 16838 22652 16890
rect 22356 16836 22412 16838
rect 22436 16836 22492 16838
rect 22516 16836 22572 16838
rect 22596 16836 22652 16838
rect 22356 15802 22412 15804
rect 22436 15802 22492 15804
rect 22516 15802 22572 15804
rect 22596 15802 22652 15804
rect 22356 15750 22402 15802
rect 22402 15750 22412 15802
rect 22436 15750 22466 15802
rect 22466 15750 22478 15802
rect 22478 15750 22492 15802
rect 22516 15750 22530 15802
rect 22530 15750 22542 15802
rect 22542 15750 22572 15802
rect 22596 15750 22606 15802
rect 22606 15750 22652 15802
rect 22356 15748 22412 15750
rect 22436 15748 22492 15750
rect 22516 15748 22572 15750
rect 22596 15748 22652 15750
rect 23662 19760 23718 19816
rect 23570 19116 23572 19136
rect 23572 19116 23624 19136
rect 23624 19116 23626 19136
rect 23570 19080 23626 19116
rect 23294 17720 23350 17776
rect 23386 16496 23442 16552
rect 23856 19610 23912 19612
rect 23936 19610 23992 19612
rect 24016 19610 24072 19612
rect 24096 19610 24152 19612
rect 23856 19558 23902 19610
rect 23902 19558 23912 19610
rect 23936 19558 23966 19610
rect 23966 19558 23978 19610
rect 23978 19558 23992 19610
rect 24016 19558 24030 19610
rect 24030 19558 24042 19610
rect 24042 19558 24072 19610
rect 24096 19558 24106 19610
rect 24106 19558 24152 19610
rect 23856 19556 23912 19558
rect 23936 19556 23992 19558
rect 24016 19556 24072 19558
rect 24096 19556 24152 19558
rect 23856 18522 23912 18524
rect 23936 18522 23992 18524
rect 24016 18522 24072 18524
rect 24096 18522 24152 18524
rect 23856 18470 23902 18522
rect 23902 18470 23912 18522
rect 23936 18470 23966 18522
rect 23966 18470 23978 18522
rect 23978 18470 23992 18522
rect 24016 18470 24030 18522
rect 24030 18470 24042 18522
rect 24042 18470 24072 18522
rect 24096 18470 24106 18522
rect 24106 18470 24152 18522
rect 23856 18468 23912 18470
rect 23936 18468 23992 18470
rect 24016 18468 24072 18470
rect 24096 18468 24152 18470
rect 24306 18400 24362 18456
rect 23856 17434 23912 17436
rect 23936 17434 23992 17436
rect 24016 17434 24072 17436
rect 24096 17434 24152 17436
rect 23856 17382 23902 17434
rect 23902 17382 23912 17434
rect 23936 17382 23966 17434
rect 23966 17382 23978 17434
rect 23978 17382 23992 17434
rect 24016 17382 24030 17434
rect 24030 17382 24042 17434
rect 24042 17382 24072 17434
rect 24096 17382 24106 17434
rect 24106 17382 24152 17434
rect 23856 17380 23912 17382
rect 23936 17380 23992 17382
rect 24016 17380 24072 17382
rect 24096 17380 24152 17382
rect 23754 17040 23810 17096
rect 23856 16346 23912 16348
rect 23936 16346 23992 16348
rect 24016 16346 24072 16348
rect 24096 16346 24152 16348
rect 23856 16294 23902 16346
rect 23902 16294 23912 16346
rect 23936 16294 23966 16346
rect 23966 16294 23978 16346
rect 23978 16294 23992 16346
rect 24016 16294 24030 16346
rect 24030 16294 24042 16346
rect 24042 16294 24072 16346
rect 24096 16294 24106 16346
rect 24106 16294 24152 16346
rect 23856 16292 23912 16294
rect 23936 16292 23992 16294
rect 24016 16292 24072 16294
rect 24096 16292 24152 16294
rect 23386 15680 23442 15736
rect 22282 15580 22284 15600
rect 22284 15580 22336 15600
rect 22336 15580 22338 15600
rect 22282 15544 22338 15580
rect 20856 11994 20912 11996
rect 20936 11994 20992 11996
rect 21016 11994 21072 11996
rect 21096 11994 21152 11996
rect 20856 11942 20902 11994
rect 20902 11942 20912 11994
rect 20936 11942 20966 11994
rect 20966 11942 20978 11994
rect 20978 11942 20992 11994
rect 21016 11942 21030 11994
rect 21030 11942 21042 11994
rect 21042 11942 21072 11994
rect 21096 11942 21106 11994
rect 21106 11942 21152 11994
rect 20856 11940 20912 11942
rect 20936 11940 20992 11942
rect 21016 11940 21072 11942
rect 21096 11940 21152 11942
rect 17856 10906 17912 10908
rect 17936 10906 17992 10908
rect 18016 10906 18072 10908
rect 18096 10906 18152 10908
rect 17856 10854 17902 10906
rect 17902 10854 17912 10906
rect 17936 10854 17966 10906
rect 17966 10854 17978 10906
rect 17978 10854 17992 10906
rect 18016 10854 18030 10906
rect 18030 10854 18042 10906
rect 18042 10854 18072 10906
rect 18096 10854 18106 10906
rect 18106 10854 18152 10906
rect 17856 10852 17912 10854
rect 17936 10852 17992 10854
rect 18016 10852 18072 10854
rect 18096 10852 18152 10854
rect 19356 10362 19412 10364
rect 19436 10362 19492 10364
rect 19516 10362 19572 10364
rect 19596 10362 19652 10364
rect 19356 10310 19402 10362
rect 19402 10310 19412 10362
rect 19436 10310 19466 10362
rect 19466 10310 19478 10362
rect 19478 10310 19492 10362
rect 19516 10310 19530 10362
rect 19530 10310 19542 10362
rect 19542 10310 19572 10362
rect 19596 10310 19606 10362
rect 19606 10310 19652 10362
rect 19356 10308 19412 10310
rect 19436 10308 19492 10310
rect 19516 10308 19572 10310
rect 19596 10308 19652 10310
rect 17856 9818 17912 9820
rect 17936 9818 17992 9820
rect 18016 9818 18072 9820
rect 18096 9818 18152 9820
rect 17856 9766 17902 9818
rect 17902 9766 17912 9818
rect 17936 9766 17966 9818
rect 17966 9766 17978 9818
rect 17978 9766 17992 9818
rect 18016 9766 18030 9818
rect 18030 9766 18042 9818
rect 18042 9766 18072 9818
rect 18096 9766 18106 9818
rect 18106 9766 18152 9818
rect 17856 9764 17912 9766
rect 17936 9764 17992 9766
rect 18016 9764 18072 9766
rect 18096 9764 18152 9766
rect 20856 10906 20912 10908
rect 20936 10906 20992 10908
rect 21016 10906 21072 10908
rect 21096 10906 21152 10908
rect 20856 10854 20902 10906
rect 20902 10854 20912 10906
rect 20936 10854 20966 10906
rect 20966 10854 20978 10906
rect 20978 10854 20992 10906
rect 21016 10854 21030 10906
rect 21030 10854 21042 10906
rect 21042 10854 21072 10906
rect 21096 10854 21106 10906
rect 21106 10854 21152 10906
rect 20856 10852 20912 10854
rect 20936 10852 20992 10854
rect 21016 10852 21072 10854
rect 21096 10852 21152 10854
rect 20856 9818 20912 9820
rect 20936 9818 20992 9820
rect 21016 9818 21072 9820
rect 21096 9818 21152 9820
rect 20856 9766 20902 9818
rect 20902 9766 20912 9818
rect 20936 9766 20966 9818
rect 20966 9766 20978 9818
rect 20978 9766 20992 9818
rect 21016 9766 21030 9818
rect 21030 9766 21042 9818
rect 21042 9766 21072 9818
rect 21096 9766 21106 9818
rect 21106 9766 21152 9818
rect 20856 9764 20912 9766
rect 20936 9764 20992 9766
rect 21016 9764 21072 9766
rect 21096 9764 21152 9766
rect 15198 8200 15254 8256
rect 13356 2746 13412 2748
rect 13436 2746 13492 2748
rect 13516 2746 13572 2748
rect 13596 2746 13652 2748
rect 13356 2694 13402 2746
rect 13402 2694 13412 2746
rect 13436 2694 13466 2746
rect 13466 2694 13478 2746
rect 13478 2694 13492 2746
rect 13516 2694 13530 2746
rect 13530 2694 13542 2746
rect 13542 2694 13572 2746
rect 13596 2694 13606 2746
rect 13606 2694 13652 2746
rect 13356 2692 13412 2694
rect 13436 2692 13492 2694
rect 13516 2692 13572 2694
rect 13596 2692 13652 2694
rect 14856 7642 14912 7644
rect 14936 7642 14992 7644
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 14856 7590 14902 7642
rect 14902 7590 14912 7642
rect 14936 7590 14966 7642
rect 14966 7590 14978 7642
rect 14978 7590 14992 7642
rect 15016 7590 15030 7642
rect 15030 7590 15042 7642
rect 15042 7590 15072 7642
rect 15096 7590 15106 7642
rect 15106 7590 15152 7642
rect 14856 7588 14912 7590
rect 14936 7588 14992 7590
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 16356 8186 16412 8188
rect 16436 8186 16492 8188
rect 16516 8186 16572 8188
rect 16596 8186 16652 8188
rect 16356 8134 16402 8186
rect 16402 8134 16412 8186
rect 16436 8134 16466 8186
rect 16466 8134 16478 8186
rect 16478 8134 16492 8186
rect 16516 8134 16530 8186
rect 16530 8134 16542 8186
rect 16542 8134 16572 8186
rect 16596 8134 16606 8186
rect 16606 8134 16652 8186
rect 16356 8132 16412 8134
rect 16436 8132 16492 8134
rect 16516 8132 16572 8134
rect 16596 8132 16652 8134
rect 17856 8730 17912 8732
rect 17936 8730 17992 8732
rect 18016 8730 18072 8732
rect 18096 8730 18152 8732
rect 17856 8678 17902 8730
rect 17902 8678 17912 8730
rect 17936 8678 17966 8730
rect 17966 8678 17978 8730
rect 17978 8678 17992 8730
rect 18016 8678 18030 8730
rect 18030 8678 18042 8730
rect 18042 8678 18072 8730
rect 18096 8678 18106 8730
rect 18106 8678 18152 8730
rect 17856 8676 17912 8678
rect 17936 8676 17992 8678
rect 18016 8676 18072 8678
rect 18096 8676 18152 8678
rect 14856 6554 14912 6556
rect 14936 6554 14992 6556
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 14856 6502 14902 6554
rect 14902 6502 14912 6554
rect 14936 6502 14966 6554
rect 14966 6502 14978 6554
rect 14978 6502 14992 6554
rect 15016 6502 15030 6554
rect 15030 6502 15042 6554
rect 15042 6502 15072 6554
rect 15096 6502 15106 6554
rect 15106 6502 15152 6554
rect 14856 6500 14912 6502
rect 14936 6500 14992 6502
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 14856 5466 14912 5468
rect 14936 5466 14992 5468
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 14856 5414 14902 5466
rect 14902 5414 14912 5466
rect 14936 5414 14966 5466
rect 14966 5414 14978 5466
rect 14978 5414 14992 5466
rect 15016 5414 15030 5466
rect 15030 5414 15042 5466
rect 15042 5414 15072 5466
rect 15096 5414 15106 5466
rect 15106 5414 15152 5466
rect 14856 5412 14912 5414
rect 14936 5412 14992 5414
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 14856 4378 14912 4380
rect 14936 4378 14992 4380
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 14856 4326 14902 4378
rect 14902 4326 14912 4378
rect 14936 4326 14966 4378
rect 14966 4326 14978 4378
rect 14978 4326 14992 4378
rect 15016 4326 15030 4378
rect 15030 4326 15042 4378
rect 15042 4326 15072 4378
rect 15096 4326 15106 4378
rect 15106 4326 15152 4378
rect 14856 4324 14912 4326
rect 14936 4324 14992 4326
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 14738 3440 14794 3496
rect 14856 3290 14912 3292
rect 14936 3290 14992 3292
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 14856 3238 14902 3290
rect 14902 3238 14912 3290
rect 14936 3238 14966 3290
rect 14966 3238 14978 3290
rect 14978 3238 14992 3290
rect 15016 3238 15030 3290
rect 15030 3238 15042 3290
rect 15042 3238 15072 3290
rect 15096 3238 15106 3290
rect 15106 3238 15152 3290
rect 14856 3236 14912 3238
rect 14936 3236 14992 3238
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 16356 7098 16412 7100
rect 16436 7098 16492 7100
rect 16516 7098 16572 7100
rect 16596 7098 16652 7100
rect 16356 7046 16402 7098
rect 16402 7046 16412 7098
rect 16436 7046 16466 7098
rect 16466 7046 16478 7098
rect 16478 7046 16492 7098
rect 16516 7046 16530 7098
rect 16530 7046 16542 7098
rect 16542 7046 16572 7098
rect 16596 7046 16606 7098
rect 16606 7046 16652 7098
rect 16356 7044 16412 7046
rect 16436 7044 16492 7046
rect 16516 7044 16572 7046
rect 16596 7044 16652 7046
rect 16356 6010 16412 6012
rect 16436 6010 16492 6012
rect 16516 6010 16572 6012
rect 16596 6010 16652 6012
rect 16356 5958 16402 6010
rect 16402 5958 16412 6010
rect 16436 5958 16466 6010
rect 16466 5958 16478 6010
rect 16478 5958 16492 6010
rect 16516 5958 16530 6010
rect 16530 5958 16542 6010
rect 16542 5958 16572 6010
rect 16596 5958 16606 6010
rect 16606 5958 16652 6010
rect 16356 5956 16412 5958
rect 16436 5956 16492 5958
rect 16516 5956 16572 5958
rect 16596 5956 16652 5958
rect 16356 4922 16412 4924
rect 16436 4922 16492 4924
rect 16516 4922 16572 4924
rect 16596 4922 16652 4924
rect 16356 4870 16402 4922
rect 16402 4870 16412 4922
rect 16436 4870 16466 4922
rect 16466 4870 16478 4922
rect 16478 4870 16492 4922
rect 16516 4870 16530 4922
rect 16530 4870 16542 4922
rect 16542 4870 16572 4922
rect 16596 4870 16606 4922
rect 16606 4870 16652 4922
rect 16356 4868 16412 4870
rect 16436 4868 16492 4870
rect 16516 4868 16572 4870
rect 16596 4868 16652 4870
rect 16356 3834 16412 3836
rect 16436 3834 16492 3836
rect 16516 3834 16572 3836
rect 16596 3834 16652 3836
rect 16356 3782 16402 3834
rect 16402 3782 16412 3834
rect 16436 3782 16466 3834
rect 16466 3782 16478 3834
rect 16478 3782 16492 3834
rect 16516 3782 16530 3834
rect 16530 3782 16542 3834
rect 16542 3782 16572 3834
rect 16596 3782 16606 3834
rect 16606 3782 16652 3834
rect 16356 3780 16412 3782
rect 16436 3780 16492 3782
rect 16516 3780 16572 3782
rect 16596 3780 16652 3782
rect 16210 3476 16212 3496
rect 16212 3476 16264 3496
rect 16264 3476 16266 3496
rect 16210 3440 16266 3476
rect 16356 2746 16412 2748
rect 16436 2746 16492 2748
rect 16516 2746 16572 2748
rect 16596 2746 16652 2748
rect 16356 2694 16402 2746
rect 16402 2694 16412 2746
rect 16436 2694 16466 2746
rect 16466 2694 16478 2746
rect 16478 2694 16492 2746
rect 16516 2694 16530 2746
rect 16530 2694 16542 2746
rect 16542 2694 16572 2746
rect 16596 2694 16606 2746
rect 16606 2694 16652 2746
rect 16356 2692 16412 2694
rect 16436 2692 16492 2694
rect 16516 2692 16572 2694
rect 16596 2692 16652 2694
rect 19356 9274 19412 9276
rect 19436 9274 19492 9276
rect 19516 9274 19572 9276
rect 19596 9274 19652 9276
rect 19356 9222 19402 9274
rect 19402 9222 19412 9274
rect 19436 9222 19466 9274
rect 19466 9222 19478 9274
rect 19478 9222 19492 9274
rect 19516 9222 19530 9274
rect 19530 9222 19542 9274
rect 19542 9222 19572 9274
rect 19596 9222 19606 9274
rect 19606 9222 19652 9274
rect 19356 9220 19412 9222
rect 19436 9220 19492 9222
rect 19516 9220 19572 9222
rect 19596 9220 19652 9222
rect 22098 13676 22100 13696
rect 22100 13676 22152 13696
rect 22152 13676 22154 13696
rect 22098 13640 22154 13676
rect 22356 14714 22412 14716
rect 22436 14714 22492 14716
rect 22516 14714 22572 14716
rect 22596 14714 22652 14716
rect 22356 14662 22402 14714
rect 22402 14662 22412 14714
rect 22436 14662 22466 14714
rect 22466 14662 22478 14714
rect 22478 14662 22492 14714
rect 22516 14662 22530 14714
rect 22530 14662 22542 14714
rect 22542 14662 22572 14714
rect 22596 14662 22606 14714
rect 22606 14662 22652 14714
rect 22356 14660 22412 14662
rect 22436 14660 22492 14662
rect 22516 14660 22572 14662
rect 22596 14660 22652 14662
rect 22356 13626 22412 13628
rect 22436 13626 22492 13628
rect 22516 13626 22572 13628
rect 22596 13626 22652 13628
rect 22356 13574 22402 13626
rect 22402 13574 22412 13626
rect 22436 13574 22466 13626
rect 22466 13574 22478 13626
rect 22478 13574 22492 13626
rect 22516 13574 22530 13626
rect 22530 13574 22542 13626
rect 22542 13574 22572 13626
rect 22596 13574 22606 13626
rect 22606 13574 22652 13626
rect 22356 13572 22412 13574
rect 22436 13572 22492 13574
rect 22516 13572 22572 13574
rect 22596 13572 22652 13574
rect 22356 12538 22412 12540
rect 22436 12538 22492 12540
rect 22516 12538 22572 12540
rect 22596 12538 22652 12540
rect 22356 12486 22402 12538
rect 22402 12486 22412 12538
rect 22436 12486 22466 12538
rect 22466 12486 22478 12538
rect 22478 12486 22492 12538
rect 22516 12486 22530 12538
rect 22530 12486 22542 12538
rect 22542 12486 22572 12538
rect 22596 12486 22606 12538
rect 22606 12486 22652 12538
rect 22356 12484 22412 12486
rect 22436 12484 22492 12486
rect 22516 12484 22572 12486
rect 22596 12484 22652 12486
rect 23856 15258 23912 15260
rect 23936 15258 23992 15260
rect 24016 15258 24072 15260
rect 24096 15258 24152 15260
rect 23856 15206 23902 15258
rect 23902 15206 23912 15258
rect 23936 15206 23966 15258
rect 23966 15206 23978 15258
rect 23978 15206 23992 15258
rect 24016 15206 24030 15258
rect 24030 15206 24042 15258
rect 24042 15206 24072 15258
rect 24096 15206 24106 15258
rect 24106 15206 24152 15258
rect 23856 15204 23912 15206
rect 23936 15204 23992 15206
rect 24016 15204 24072 15206
rect 24096 15204 24152 15206
rect 23570 14320 23626 14376
rect 23856 14170 23912 14172
rect 23936 14170 23992 14172
rect 24016 14170 24072 14172
rect 24096 14170 24152 14172
rect 23856 14118 23902 14170
rect 23902 14118 23912 14170
rect 23936 14118 23966 14170
rect 23966 14118 23978 14170
rect 23978 14118 23992 14170
rect 24016 14118 24030 14170
rect 24030 14118 24042 14170
rect 24042 14118 24072 14170
rect 24096 14118 24106 14170
rect 24106 14118 24152 14170
rect 23856 14116 23912 14118
rect 23936 14116 23992 14118
rect 24016 14116 24072 14118
rect 24096 14116 24152 14118
rect 23662 13640 23718 13696
rect 22356 11450 22412 11452
rect 22436 11450 22492 11452
rect 22516 11450 22572 11452
rect 22596 11450 22652 11452
rect 22356 11398 22402 11450
rect 22402 11398 22412 11450
rect 22436 11398 22466 11450
rect 22466 11398 22478 11450
rect 22478 11398 22492 11450
rect 22516 11398 22530 11450
rect 22530 11398 22542 11450
rect 22542 11398 22572 11450
rect 22596 11398 22606 11450
rect 22606 11398 22652 11450
rect 22356 11396 22412 11398
rect 22436 11396 22492 11398
rect 22516 11396 22572 11398
rect 22596 11396 22652 11398
rect 19356 8186 19412 8188
rect 19436 8186 19492 8188
rect 19516 8186 19572 8188
rect 19596 8186 19652 8188
rect 19356 8134 19402 8186
rect 19402 8134 19412 8186
rect 19436 8134 19466 8186
rect 19466 8134 19478 8186
rect 19478 8134 19492 8186
rect 19516 8134 19530 8186
rect 19530 8134 19542 8186
rect 19542 8134 19572 8186
rect 19596 8134 19606 8186
rect 19606 8134 19652 8186
rect 19356 8132 19412 8134
rect 19436 8132 19492 8134
rect 19516 8132 19572 8134
rect 19596 8132 19652 8134
rect 17856 7642 17912 7644
rect 17936 7642 17992 7644
rect 18016 7642 18072 7644
rect 18096 7642 18152 7644
rect 17856 7590 17902 7642
rect 17902 7590 17912 7642
rect 17936 7590 17966 7642
rect 17966 7590 17978 7642
rect 17978 7590 17992 7642
rect 18016 7590 18030 7642
rect 18030 7590 18042 7642
rect 18042 7590 18072 7642
rect 18096 7590 18106 7642
rect 18106 7590 18152 7642
rect 17856 7588 17912 7590
rect 17936 7588 17992 7590
rect 18016 7588 18072 7590
rect 18096 7588 18152 7590
rect 17856 6554 17912 6556
rect 17936 6554 17992 6556
rect 18016 6554 18072 6556
rect 18096 6554 18152 6556
rect 17856 6502 17902 6554
rect 17902 6502 17912 6554
rect 17936 6502 17966 6554
rect 17966 6502 17978 6554
rect 17978 6502 17992 6554
rect 18016 6502 18030 6554
rect 18030 6502 18042 6554
rect 18042 6502 18072 6554
rect 18096 6502 18106 6554
rect 18106 6502 18152 6554
rect 17856 6500 17912 6502
rect 17936 6500 17992 6502
rect 18016 6500 18072 6502
rect 18096 6500 18152 6502
rect 17856 5466 17912 5468
rect 17936 5466 17992 5468
rect 18016 5466 18072 5468
rect 18096 5466 18152 5468
rect 17856 5414 17902 5466
rect 17902 5414 17912 5466
rect 17936 5414 17966 5466
rect 17966 5414 17978 5466
rect 17978 5414 17992 5466
rect 18016 5414 18030 5466
rect 18030 5414 18042 5466
rect 18042 5414 18072 5466
rect 18096 5414 18106 5466
rect 18106 5414 18152 5466
rect 17856 5412 17912 5414
rect 17936 5412 17992 5414
rect 18016 5412 18072 5414
rect 18096 5412 18152 5414
rect 17856 4378 17912 4380
rect 17936 4378 17992 4380
rect 18016 4378 18072 4380
rect 18096 4378 18152 4380
rect 17856 4326 17902 4378
rect 17902 4326 17912 4378
rect 17936 4326 17966 4378
rect 17966 4326 17978 4378
rect 17978 4326 17992 4378
rect 18016 4326 18030 4378
rect 18030 4326 18042 4378
rect 18042 4326 18072 4378
rect 18096 4326 18106 4378
rect 18106 4326 18152 4378
rect 17856 4324 17912 4326
rect 17936 4324 17992 4326
rect 18016 4324 18072 4326
rect 18096 4324 18152 4326
rect 17856 3290 17912 3292
rect 17936 3290 17992 3292
rect 18016 3290 18072 3292
rect 18096 3290 18152 3292
rect 17856 3238 17902 3290
rect 17902 3238 17912 3290
rect 17936 3238 17966 3290
rect 17966 3238 17978 3290
rect 17978 3238 17992 3290
rect 18016 3238 18030 3290
rect 18030 3238 18042 3290
rect 18042 3238 18072 3290
rect 18096 3238 18106 3290
rect 18106 3238 18152 3290
rect 17856 3236 17912 3238
rect 17936 3236 17992 3238
rect 18016 3236 18072 3238
rect 18096 3236 18152 3238
rect 2856 2202 2912 2204
rect 2936 2202 2992 2204
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 2856 2150 2902 2202
rect 2902 2150 2912 2202
rect 2936 2150 2966 2202
rect 2966 2150 2978 2202
rect 2978 2150 2992 2202
rect 3016 2150 3030 2202
rect 3030 2150 3042 2202
rect 3042 2150 3072 2202
rect 3096 2150 3106 2202
rect 3106 2150 3152 2202
rect 2856 2148 2912 2150
rect 2936 2148 2992 2150
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 5856 2202 5912 2204
rect 5936 2202 5992 2204
rect 6016 2202 6072 2204
rect 6096 2202 6152 2204
rect 5856 2150 5902 2202
rect 5902 2150 5912 2202
rect 5936 2150 5966 2202
rect 5966 2150 5978 2202
rect 5978 2150 5992 2202
rect 6016 2150 6030 2202
rect 6030 2150 6042 2202
rect 6042 2150 6072 2202
rect 6096 2150 6106 2202
rect 6106 2150 6152 2202
rect 5856 2148 5912 2150
rect 5936 2148 5992 2150
rect 6016 2148 6072 2150
rect 6096 2148 6152 2150
rect 8856 2202 8912 2204
rect 8936 2202 8992 2204
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 8856 2150 8902 2202
rect 8902 2150 8912 2202
rect 8936 2150 8966 2202
rect 8966 2150 8978 2202
rect 8978 2150 8992 2202
rect 9016 2150 9030 2202
rect 9030 2150 9042 2202
rect 9042 2150 9072 2202
rect 9096 2150 9106 2202
rect 9106 2150 9152 2202
rect 8856 2148 8912 2150
rect 8936 2148 8992 2150
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 11856 2202 11912 2204
rect 11936 2202 11992 2204
rect 12016 2202 12072 2204
rect 12096 2202 12152 2204
rect 11856 2150 11902 2202
rect 11902 2150 11912 2202
rect 11936 2150 11966 2202
rect 11966 2150 11978 2202
rect 11978 2150 11992 2202
rect 12016 2150 12030 2202
rect 12030 2150 12042 2202
rect 12042 2150 12072 2202
rect 12096 2150 12106 2202
rect 12106 2150 12152 2202
rect 11856 2148 11912 2150
rect 11936 2148 11992 2150
rect 12016 2148 12072 2150
rect 12096 2148 12152 2150
rect 14856 2202 14912 2204
rect 14936 2202 14992 2204
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 14856 2150 14902 2202
rect 14902 2150 14912 2202
rect 14936 2150 14966 2202
rect 14966 2150 14978 2202
rect 14978 2150 14992 2202
rect 15016 2150 15030 2202
rect 15030 2150 15042 2202
rect 15042 2150 15072 2202
rect 15096 2150 15106 2202
rect 15106 2150 15152 2202
rect 14856 2148 14912 2150
rect 14936 2148 14992 2150
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 19356 7098 19412 7100
rect 19436 7098 19492 7100
rect 19516 7098 19572 7100
rect 19596 7098 19652 7100
rect 19356 7046 19402 7098
rect 19402 7046 19412 7098
rect 19436 7046 19466 7098
rect 19466 7046 19478 7098
rect 19478 7046 19492 7098
rect 19516 7046 19530 7098
rect 19530 7046 19542 7098
rect 19542 7046 19572 7098
rect 19596 7046 19606 7098
rect 19606 7046 19652 7098
rect 19356 7044 19412 7046
rect 19436 7044 19492 7046
rect 19516 7044 19572 7046
rect 19596 7044 19652 7046
rect 19356 6010 19412 6012
rect 19436 6010 19492 6012
rect 19516 6010 19572 6012
rect 19596 6010 19652 6012
rect 19356 5958 19402 6010
rect 19402 5958 19412 6010
rect 19436 5958 19466 6010
rect 19466 5958 19478 6010
rect 19478 5958 19492 6010
rect 19516 5958 19530 6010
rect 19530 5958 19542 6010
rect 19542 5958 19572 6010
rect 19596 5958 19606 6010
rect 19606 5958 19652 6010
rect 19356 5956 19412 5958
rect 19436 5956 19492 5958
rect 19516 5956 19572 5958
rect 19596 5956 19652 5958
rect 19356 4922 19412 4924
rect 19436 4922 19492 4924
rect 19516 4922 19572 4924
rect 19596 4922 19652 4924
rect 19356 4870 19402 4922
rect 19402 4870 19412 4922
rect 19436 4870 19466 4922
rect 19466 4870 19478 4922
rect 19478 4870 19492 4922
rect 19516 4870 19530 4922
rect 19530 4870 19542 4922
rect 19542 4870 19572 4922
rect 19596 4870 19606 4922
rect 19606 4870 19652 4922
rect 19356 4868 19412 4870
rect 19436 4868 19492 4870
rect 19516 4868 19572 4870
rect 19596 4868 19652 4870
rect 19356 3834 19412 3836
rect 19436 3834 19492 3836
rect 19516 3834 19572 3836
rect 19596 3834 19652 3836
rect 19356 3782 19402 3834
rect 19402 3782 19412 3834
rect 19436 3782 19466 3834
rect 19466 3782 19478 3834
rect 19478 3782 19492 3834
rect 19516 3782 19530 3834
rect 19530 3782 19542 3834
rect 19542 3782 19572 3834
rect 19596 3782 19606 3834
rect 19606 3782 19652 3834
rect 19356 3780 19412 3782
rect 19436 3780 19492 3782
rect 19516 3780 19572 3782
rect 19596 3780 19652 3782
rect 20856 8730 20912 8732
rect 20936 8730 20992 8732
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 20856 8678 20902 8730
rect 20902 8678 20912 8730
rect 20936 8678 20966 8730
rect 20966 8678 20978 8730
rect 20978 8678 20992 8730
rect 21016 8678 21030 8730
rect 21030 8678 21042 8730
rect 21042 8678 21072 8730
rect 21096 8678 21106 8730
rect 21106 8678 21152 8730
rect 20856 8676 20912 8678
rect 20936 8676 20992 8678
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 20626 8336 20682 8392
rect 20856 7642 20912 7644
rect 20936 7642 20992 7644
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 20856 7590 20902 7642
rect 20902 7590 20912 7642
rect 20936 7590 20966 7642
rect 20966 7590 20978 7642
rect 20978 7590 20992 7642
rect 21016 7590 21030 7642
rect 21030 7590 21042 7642
rect 21042 7590 21072 7642
rect 21096 7590 21106 7642
rect 21106 7590 21152 7642
rect 20856 7588 20912 7590
rect 20936 7588 20992 7590
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 20856 6554 20912 6556
rect 20936 6554 20992 6556
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 20856 6502 20902 6554
rect 20902 6502 20912 6554
rect 20936 6502 20966 6554
rect 20966 6502 20978 6554
rect 20978 6502 20992 6554
rect 21016 6502 21030 6554
rect 21030 6502 21042 6554
rect 21042 6502 21072 6554
rect 21096 6502 21106 6554
rect 21106 6502 21152 6554
rect 20856 6500 20912 6502
rect 20936 6500 20992 6502
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 22356 10362 22412 10364
rect 22436 10362 22492 10364
rect 22516 10362 22572 10364
rect 22596 10362 22652 10364
rect 22356 10310 22402 10362
rect 22402 10310 22412 10362
rect 22436 10310 22466 10362
rect 22466 10310 22478 10362
rect 22478 10310 22492 10362
rect 22516 10310 22530 10362
rect 22530 10310 22542 10362
rect 22542 10310 22572 10362
rect 22596 10310 22606 10362
rect 22606 10310 22652 10362
rect 22356 10308 22412 10310
rect 22436 10308 22492 10310
rect 22516 10308 22572 10310
rect 22596 10308 22652 10310
rect 23570 12316 23572 12336
rect 23572 12316 23624 12336
rect 23624 12316 23626 12336
rect 23570 12280 23626 12316
rect 23856 13082 23912 13084
rect 23936 13082 23992 13084
rect 24016 13082 24072 13084
rect 24096 13082 24152 13084
rect 23856 13030 23902 13082
rect 23902 13030 23912 13082
rect 23936 13030 23966 13082
rect 23966 13030 23978 13082
rect 23978 13030 23992 13082
rect 24016 13030 24030 13082
rect 24030 13030 24042 13082
rect 24042 13030 24072 13082
rect 24096 13030 24106 13082
rect 24106 13030 24152 13082
rect 23856 13028 23912 13030
rect 23936 13028 23992 13030
rect 24016 13028 24072 13030
rect 24096 13028 24152 13030
rect 24306 12960 24362 13016
rect 23856 11994 23912 11996
rect 23936 11994 23992 11996
rect 24016 11994 24072 11996
rect 24096 11994 24152 11996
rect 23856 11942 23902 11994
rect 23902 11942 23912 11994
rect 23936 11942 23966 11994
rect 23966 11942 23978 11994
rect 23978 11942 23992 11994
rect 24016 11942 24030 11994
rect 24030 11942 24042 11994
rect 24042 11942 24072 11994
rect 24096 11942 24106 11994
rect 24106 11942 24152 11994
rect 23856 11940 23912 11942
rect 23936 11940 23992 11942
rect 24016 11940 24072 11942
rect 24096 11940 24152 11942
rect 23478 11600 23534 11656
rect 23856 10906 23912 10908
rect 23936 10906 23992 10908
rect 24016 10906 24072 10908
rect 24096 10906 24152 10908
rect 23856 10854 23902 10906
rect 23902 10854 23912 10906
rect 23936 10854 23966 10906
rect 23966 10854 23978 10906
rect 23978 10854 23992 10906
rect 24016 10854 24030 10906
rect 24030 10854 24042 10906
rect 24042 10854 24072 10906
rect 24096 10854 24106 10906
rect 24106 10854 24152 10906
rect 23856 10852 23912 10854
rect 23936 10852 23992 10854
rect 24016 10852 24072 10854
rect 24096 10852 24152 10854
rect 23294 10648 23350 10704
rect 22356 9274 22412 9276
rect 22436 9274 22492 9276
rect 22516 9274 22572 9276
rect 22596 9274 22652 9276
rect 22356 9222 22402 9274
rect 22402 9222 22412 9274
rect 22436 9222 22466 9274
rect 22466 9222 22478 9274
rect 22478 9222 22492 9274
rect 22516 9222 22530 9274
rect 22530 9222 22542 9274
rect 22542 9222 22572 9274
rect 22596 9222 22606 9274
rect 22606 9222 22652 9274
rect 22356 9220 22412 9222
rect 22436 9220 22492 9222
rect 22516 9220 22572 9222
rect 22596 9220 22652 9222
rect 22834 9560 22890 9616
rect 23386 10240 23442 10296
rect 23856 9818 23912 9820
rect 23936 9818 23992 9820
rect 24016 9818 24072 9820
rect 24096 9818 24152 9820
rect 23856 9766 23902 9818
rect 23902 9766 23912 9818
rect 23936 9766 23966 9818
rect 23966 9766 23978 9818
rect 23978 9766 23992 9818
rect 24016 9766 24030 9818
rect 24030 9766 24042 9818
rect 24042 9766 24072 9818
rect 24096 9766 24106 9818
rect 24106 9766 24152 9818
rect 23856 9764 23912 9766
rect 23936 9764 23992 9766
rect 24016 9764 24072 9766
rect 24096 9764 24152 9766
rect 23386 8916 23388 8936
rect 23388 8916 23440 8936
rect 23440 8916 23442 8936
rect 23386 8880 23442 8916
rect 23856 8730 23912 8732
rect 23936 8730 23992 8732
rect 24016 8730 24072 8732
rect 24096 8730 24152 8732
rect 23856 8678 23902 8730
rect 23902 8678 23912 8730
rect 23936 8678 23966 8730
rect 23966 8678 23978 8730
rect 23978 8678 23992 8730
rect 24016 8678 24030 8730
rect 24030 8678 24042 8730
rect 24042 8678 24072 8730
rect 24096 8678 24106 8730
rect 24106 8678 24152 8730
rect 23856 8676 23912 8678
rect 23936 8676 23992 8678
rect 24016 8676 24072 8678
rect 24096 8676 24152 8678
rect 22356 8186 22412 8188
rect 22436 8186 22492 8188
rect 22516 8186 22572 8188
rect 22596 8186 22652 8188
rect 22356 8134 22402 8186
rect 22402 8134 22412 8186
rect 22436 8134 22466 8186
rect 22466 8134 22478 8186
rect 22478 8134 22492 8186
rect 22516 8134 22530 8186
rect 22530 8134 22542 8186
rect 22542 8134 22572 8186
rect 22596 8134 22606 8186
rect 22606 8134 22652 8186
rect 22356 8132 22412 8134
rect 22436 8132 22492 8134
rect 22516 8132 22572 8134
rect 22596 8132 22652 8134
rect 23856 7642 23912 7644
rect 23936 7642 23992 7644
rect 24016 7642 24072 7644
rect 24096 7642 24152 7644
rect 23856 7590 23902 7642
rect 23902 7590 23912 7642
rect 23936 7590 23966 7642
rect 23966 7590 23978 7642
rect 23978 7590 23992 7642
rect 24016 7590 24030 7642
rect 24030 7590 24042 7642
rect 24042 7590 24072 7642
rect 24096 7590 24106 7642
rect 24106 7590 24152 7642
rect 23856 7588 23912 7590
rect 23936 7588 23992 7590
rect 24016 7588 24072 7590
rect 24096 7588 24152 7590
rect 22356 7098 22412 7100
rect 22436 7098 22492 7100
rect 22516 7098 22572 7100
rect 22596 7098 22652 7100
rect 22356 7046 22402 7098
rect 22402 7046 22412 7098
rect 22436 7046 22466 7098
rect 22466 7046 22478 7098
rect 22478 7046 22492 7098
rect 22516 7046 22530 7098
rect 22530 7046 22542 7098
rect 22542 7046 22572 7098
rect 22596 7046 22606 7098
rect 22606 7046 22652 7098
rect 22356 7044 22412 7046
rect 22436 7044 22492 7046
rect 22516 7044 22572 7046
rect 22596 7044 22652 7046
rect 23386 6840 23442 6896
rect 23856 6554 23912 6556
rect 23936 6554 23992 6556
rect 24016 6554 24072 6556
rect 24096 6554 24152 6556
rect 23856 6502 23902 6554
rect 23902 6502 23912 6554
rect 23936 6502 23966 6554
rect 23966 6502 23978 6554
rect 23978 6502 23992 6554
rect 24016 6502 24030 6554
rect 24030 6502 24042 6554
rect 24042 6502 24072 6554
rect 24096 6502 24106 6554
rect 24106 6502 24152 6554
rect 23856 6500 23912 6502
rect 23936 6500 23992 6502
rect 24016 6500 24072 6502
rect 24096 6500 24152 6502
rect 23662 6160 23718 6216
rect 22356 6010 22412 6012
rect 22436 6010 22492 6012
rect 22516 6010 22572 6012
rect 22596 6010 22652 6012
rect 22356 5958 22402 6010
rect 22402 5958 22412 6010
rect 22436 5958 22466 6010
rect 22466 5958 22478 6010
rect 22478 5958 22492 6010
rect 22516 5958 22530 6010
rect 22530 5958 22542 6010
rect 22542 5958 22572 6010
rect 22596 5958 22606 6010
rect 22606 5958 22652 6010
rect 22356 5956 22412 5958
rect 22436 5956 22492 5958
rect 22516 5956 22572 5958
rect 22596 5956 22652 5958
rect 20856 5466 20912 5468
rect 20936 5466 20992 5468
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 20856 5414 20902 5466
rect 20902 5414 20912 5466
rect 20936 5414 20966 5466
rect 20966 5414 20978 5466
rect 20978 5414 20992 5466
rect 21016 5414 21030 5466
rect 21030 5414 21042 5466
rect 21042 5414 21072 5466
rect 21096 5414 21106 5466
rect 21106 5414 21152 5466
rect 20856 5412 20912 5414
rect 20936 5412 20992 5414
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 23856 5466 23912 5468
rect 23936 5466 23992 5468
rect 24016 5466 24072 5468
rect 24096 5466 24152 5468
rect 23856 5414 23902 5466
rect 23902 5414 23912 5466
rect 23936 5414 23966 5466
rect 23966 5414 23978 5466
rect 23978 5414 23992 5466
rect 24016 5414 24030 5466
rect 24030 5414 24042 5466
rect 24042 5414 24072 5466
rect 24096 5414 24106 5466
rect 24106 5414 24152 5466
rect 23856 5412 23912 5414
rect 23936 5412 23992 5414
rect 24016 5412 24072 5414
rect 24096 5412 24152 5414
rect 20856 4378 20912 4380
rect 20936 4378 20992 4380
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 20856 4326 20902 4378
rect 20902 4326 20912 4378
rect 20936 4326 20966 4378
rect 20966 4326 20978 4378
rect 20978 4326 20992 4378
rect 21016 4326 21030 4378
rect 21030 4326 21042 4378
rect 21042 4326 21072 4378
rect 21096 4326 21106 4378
rect 21106 4326 21152 4378
rect 20856 4324 20912 4326
rect 20936 4324 20992 4326
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 20856 3290 20912 3292
rect 20936 3290 20992 3292
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 20856 3238 20902 3290
rect 20902 3238 20912 3290
rect 20936 3238 20966 3290
rect 20966 3238 20978 3290
rect 20978 3238 20992 3290
rect 21016 3238 21030 3290
rect 21030 3238 21042 3290
rect 21042 3238 21072 3290
rect 21096 3238 21106 3290
rect 21106 3238 21152 3290
rect 20856 3236 20912 3238
rect 20936 3236 20992 3238
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 22356 4922 22412 4924
rect 22436 4922 22492 4924
rect 22516 4922 22572 4924
rect 22596 4922 22652 4924
rect 22356 4870 22402 4922
rect 22402 4870 22412 4922
rect 22436 4870 22466 4922
rect 22466 4870 22478 4922
rect 22478 4870 22492 4922
rect 22516 4870 22530 4922
rect 22530 4870 22542 4922
rect 22542 4870 22572 4922
rect 22596 4870 22606 4922
rect 22606 4870 22652 4922
rect 22356 4868 22412 4870
rect 22436 4868 22492 4870
rect 22516 4868 22572 4870
rect 22596 4868 22652 4870
rect 23856 4378 23912 4380
rect 23936 4378 23992 4380
rect 24016 4378 24072 4380
rect 24096 4378 24152 4380
rect 23856 4326 23902 4378
rect 23902 4326 23912 4378
rect 23936 4326 23966 4378
rect 23966 4326 23978 4378
rect 23978 4326 23992 4378
rect 24016 4326 24030 4378
rect 24030 4326 24042 4378
rect 24042 4326 24072 4378
rect 24096 4326 24106 4378
rect 24106 4326 24152 4378
rect 23856 4324 23912 4326
rect 23936 4324 23992 4326
rect 24016 4324 24072 4326
rect 24096 4324 24152 4326
rect 22356 3834 22412 3836
rect 22436 3834 22492 3836
rect 22516 3834 22572 3836
rect 22596 3834 22652 3836
rect 22356 3782 22402 3834
rect 22402 3782 22412 3834
rect 22436 3782 22466 3834
rect 22466 3782 22478 3834
rect 22478 3782 22492 3834
rect 22516 3782 22530 3834
rect 22530 3782 22542 3834
rect 22542 3782 22572 3834
rect 22596 3782 22606 3834
rect 22606 3782 22652 3834
rect 22356 3780 22412 3782
rect 22436 3780 22492 3782
rect 22516 3780 22572 3782
rect 22596 3780 22652 3782
rect 19356 2746 19412 2748
rect 19436 2746 19492 2748
rect 19516 2746 19572 2748
rect 19596 2746 19652 2748
rect 19356 2694 19402 2746
rect 19402 2694 19412 2746
rect 19436 2694 19466 2746
rect 19466 2694 19478 2746
rect 19478 2694 19492 2746
rect 19516 2694 19530 2746
rect 19530 2694 19542 2746
rect 19542 2694 19572 2746
rect 19596 2694 19606 2746
rect 19606 2694 19652 2746
rect 19356 2692 19412 2694
rect 19436 2692 19492 2694
rect 19516 2692 19572 2694
rect 19596 2692 19652 2694
rect 23856 3290 23912 3292
rect 23936 3290 23992 3292
rect 24016 3290 24072 3292
rect 24096 3290 24152 3292
rect 23856 3238 23902 3290
rect 23902 3238 23912 3290
rect 23936 3238 23966 3290
rect 23966 3238 23978 3290
rect 23978 3238 23992 3290
rect 24016 3238 24030 3290
rect 24030 3238 24042 3290
rect 24042 3238 24072 3290
rect 24096 3238 24106 3290
rect 24106 3238 24152 3290
rect 23856 3236 23912 3238
rect 23936 3236 23992 3238
rect 24016 3236 24072 3238
rect 24096 3236 24152 3238
rect 22356 2746 22412 2748
rect 22436 2746 22492 2748
rect 22516 2746 22572 2748
rect 22596 2746 22652 2748
rect 22356 2694 22402 2746
rect 22402 2694 22412 2746
rect 22436 2694 22466 2746
rect 22466 2694 22478 2746
rect 22478 2694 22492 2746
rect 22516 2694 22530 2746
rect 22530 2694 22542 2746
rect 22542 2694 22572 2746
rect 22596 2694 22606 2746
rect 22606 2694 22652 2746
rect 22356 2692 22412 2694
rect 22436 2692 22492 2694
rect 22516 2692 22572 2694
rect 22596 2692 22652 2694
rect 17856 2202 17912 2204
rect 17936 2202 17992 2204
rect 18016 2202 18072 2204
rect 18096 2202 18152 2204
rect 17856 2150 17902 2202
rect 17902 2150 17912 2202
rect 17936 2150 17966 2202
rect 17966 2150 17978 2202
rect 17978 2150 17992 2202
rect 18016 2150 18030 2202
rect 18030 2150 18042 2202
rect 18042 2150 18072 2202
rect 18096 2150 18106 2202
rect 18106 2150 18152 2202
rect 17856 2148 17912 2150
rect 17936 2148 17992 2150
rect 18016 2148 18072 2150
rect 18096 2148 18152 2150
rect 20856 2202 20912 2204
rect 20936 2202 20992 2204
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 20856 2150 20902 2202
rect 20902 2150 20912 2202
rect 20936 2150 20966 2202
rect 20966 2150 20978 2202
rect 20978 2150 20992 2202
rect 21016 2150 21030 2202
rect 21030 2150 21042 2202
rect 21042 2150 21072 2202
rect 21096 2150 21106 2202
rect 21106 2150 21152 2202
rect 20856 2148 20912 2150
rect 20936 2148 20992 2150
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 23856 2202 23912 2204
rect 23936 2202 23992 2204
rect 24016 2202 24072 2204
rect 24096 2202 24152 2204
rect 23856 2150 23902 2202
rect 23902 2150 23912 2202
rect 23936 2150 23966 2202
rect 23966 2150 23978 2202
rect 23978 2150 23992 2202
rect 24016 2150 24030 2202
rect 24030 2150 24042 2202
rect 24042 2150 24072 2202
rect 24096 2150 24106 2202
rect 24106 2150 24152 2202
rect 23856 2148 23912 2150
rect 23936 2148 23992 2150
rect 24016 2148 24072 2150
rect 24096 2148 24152 2150
<< metal3 >>
rect 2846 25056 3162 25057
rect 2846 24992 2852 25056
rect 2916 24992 2932 25056
rect 2996 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3162 25056
rect 2846 24991 3162 24992
rect 5846 25056 6162 25057
rect 5846 24992 5852 25056
rect 5916 24992 5932 25056
rect 5996 24992 6012 25056
rect 6076 24992 6092 25056
rect 6156 24992 6162 25056
rect 5846 24991 6162 24992
rect 8846 25056 9162 25057
rect 8846 24992 8852 25056
rect 8916 24992 8932 25056
rect 8996 24992 9012 25056
rect 9076 24992 9092 25056
rect 9156 24992 9162 25056
rect 8846 24991 9162 24992
rect 11846 25056 12162 25057
rect 11846 24992 11852 25056
rect 11916 24992 11932 25056
rect 11996 24992 12012 25056
rect 12076 24992 12092 25056
rect 12156 24992 12162 25056
rect 11846 24991 12162 24992
rect 14846 25056 15162 25057
rect 14846 24992 14852 25056
rect 14916 24992 14932 25056
rect 14996 24992 15012 25056
rect 15076 24992 15092 25056
rect 15156 24992 15162 25056
rect 14846 24991 15162 24992
rect 17846 25056 18162 25057
rect 17846 24992 17852 25056
rect 17916 24992 17932 25056
rect 17996 24992 18012 25056
rect 18076 24992 18092 25056
rect 18156 24992 18162 25056
rect 17846 24991 18162 24992
rect 20846 25056 21162 25057
rect 20846 24992 20852 25056
rect 20916 24992 20932 25056
rect 20996 24992 21012 25056
rect 21076 24992 21092 25056
rect 21156 24992 21162 25056
rect 20846 24991 21162 24992
rect 23846 25056 24162 25057
rect 23846 24992 23852 25056
rect 23916 24992 23932 25056
rect 23996 24992 24012 25056
rect 24076 24992 24092 25056
rect 24156 24992 24162 25056
rect 23846 24991 24162 24992
rect 1346 24512 1662 24513
rect 1346 24448 1352 24512
rect 1416 24448 1432 24512
rect 1496 24448 1512 24512
rect 1576 24448 1592 24512
rect 1656 24448 1662 24512
rect 1346 24447 1662 24448
rect 4346 24512 4662 24513
rect 4346 24448 4352 24512
rect 4416 24448 4432 24512
rect 4496 24448 4512 24512
rect 4576 24448 4592 24512
rect 4656 24448 4662 24512
rect 4346 24447 4662 24448
rect 7346 24512 7662 24513
rect 7346 24448 7352 24512
rect 7416 24448 7432 24512
rect 7496 24448 7512 24512
rect 7576 24448 7592 24512
rect 7656 24448 7662 24512
rect 7346 24447 7662 24448
rect 10346 24512 10662 24513
rect 10346 24448 10352 24512
rect 10416 24448 10432 24512
rect 10496 24448 10512 24512
rect 10576 24448 10592 24512
rect 10656 24448 10662 24512
rect 10346 24447 10662 24448
rect 13346 24512 13662 24513
rect 13346 24448 13352 24512
rect 13416 24448 13432 24512
rect 13496 24448 13512 24512
rect 13576 24448 13592 24512
rect 13656 24448 13662 24512
rect 13346 24447 13662 24448
rect 16346 24512 16662 24513
rect 16346 24448 16352 24512
rect 16416 24448 16432 24512
rect 16496 24448 16512 24512
rect 16576 24448 16592 24512
rect 16656 24448 16662 24512
rect 16346 24447 16662 24448
rect 19346 24512 19662 24513
rect 19346 24448 19352 24512
rect 19416 24448 19432 24512
rect 19496 24448 19512 24512
rect 19576 24448 19592 24512
rect 19656 24448 19662 24512
rect 19346 24447 19662 24448
rect 22346 24512 22662 24513
rect 22346 24448 22352 24512
rect 22416 24448 22432 24512
rect 22496 24448 22512 24512
rect 22576 24448 22592 24512
rect 22656 24448 22662 24512
rect 22346 24447 22662 24448
rect 2846 23968 3162 23969
rect 2846 23904 2852 23968
rect 2916 23904 2932 23968
rect 2996 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3162 23968
rect 2846 23903 3162 23904
rect 5846 23968 6162 23969
rect 5846 23904 5852 23968
rect 5916 23904 5932 23968
rect 5996 23904 6012 23968
rect 6076 23904 6092 23968
rect 6156 23904 6162 23968
rect 5846 23903 6162 23904
rect 8846 23968 9162 23969
rect 8846 23904 8852 23968
rect 8916 23904 8932 23968
rect 8996 23904 9012 23968
rect 9076 23904 9092 23968
rect 9156 23904 9162 23968
rect 8846 23903 9162 23904
rect 11846 23968 12162 23969
rect 11846 23904 11852 23968
rect 11916 23904 11932 23968
rect 11996 23904 12012 23968
rect 12076 23904 12092 23968
rect 12156 23904 12162 23968
rect 11846 23903 12162 23904
rect 14846 23968 15162 23969
rect 14846 23904 14852 23968
rect 14916 23904 14932 23968
rect 14996 23904 15012 23968
rect 15076 23904 15092 23968
rect 15156 23904 15162 23968
rect 14846 23903 15162 23904
rect 17846 23968 18162 23969
rect 17846 23904 17852 23968
rect 17916 23904 17932 23968
rect 17996 23904 18012 23968
rect 18076 23904 18092 23968
rect 18156 23904 18162 23968
rect 17846 23903 18162 23904
rect 20846 23968 21162 23969
rect 20846 23904 20852 23968
rect 20916 23904 20932 23968
rect 20996 23904 21012 23968
rect 21076 23904 21092 23968
rect 21156 23904 21162 23968
rect 20846 23903 21162 23904
rect 23846 23968 24162 23969
rect 23846 23904 23852 23968
rect 23916 23904 23932 23968
rect 23996 23904 24012 23968
rect 24076 23904 24092 23968
rect 24156 23904 24162 23968
rect 23846 23903 24162 23904
rect 11237 23626 11303 23629
rect 14089 23626 14155 23629
rect 15101 23626 15167 23629
rect 18781 23626 18847 23629
rect 19149 23626 19215 23629
rect 11237 23624 19215 23626
rect 11237 23568 11242 23624
rect 11298 23568 14094 23624
rect 14150 23568 15106 23624
rect 15162 23568 18786 23624
rect 18842 23568 19154 23624
rect 19210 23568 19215 23624
rect 11237 23566 19215 23568
rect 11237 23563 11303 23566
rect 14089 23563 14155 23566
rect 15101 23563 15167 23566
rect 18781 23563 18847 23566
rect 19149 23563 19215 23566
rect 1346 23424 1662 23425
rect 1346 23360 1352 23424
rect 1416 23360 1432 23424
rect 1496 23360 1512 23424
rect 1576 23360 1592 23424
rect 1656 23360 1662 23424
rect 1346 23359 1662 23360
rect 4346 23424 4662 23425
rect 4346 23360 4352 23424
rect 4416 23360 4432 23424
rect 4496 23360 4512 23424
rect 4576 23360 4592 23424
rect 4656 23360 4662 23424
rect 4346 23359 4662 23360
rect 7346 23424 7662 23425
rect 7346 23360 7352 23424
rect 7416 23360 7432 23424
rect 7496 23360 7512 23424
rect 7576 23360 7592 23424
rect 7656 23360 7662 23424
rect 7346 23359 7662 23360
rect 10346 23424 10662 23425
rect 10346 23360 10352 23424
rect 10416 23360 10432 23424
rect 10496 23360 10512 23424
rect 10576 23360 10592 23424
rect 10656 23360 10662 23424
rect 10346 23359 10662 23360
rect 13346 23424 13662 23425
rect 13346 23360 13352 23424
rect 13416 23360 13432 23424
rect 13496 23360 13512 23424
rect 13576 23360 13592 23424
rect 13656 23360 13662 23424
rect 13346 23359 13662 23360
rect 16346 23424 16662 23425
rect 16346 23360 16352 23424
rect 16416 23360 16432 23424
rect 16496 23360 16512 23424
rect 16576 23360 16592 23424
rect 16656 23360 16662 23424
rect 16346 23359 16662 23360
rect 19346 23424 19662 23425
rect 19346 23360 19352 23424
rect 19416 23360 19432 23424
rect 19496 23360 19512 23424
rect 19576 23360 19592 23424
rect 19656 23360 19662 23424
rect 19346 23359 19662 23360
rect 22346 23424 22662 23425
rect 22346 23360 22352 23424
rect 22416 23360 22432 23424
rect 22496 23360 22512 23424
rect 22576 23360 22592 23424
rect 22656 23360 22662 23424
rect 22346 23359 22662 23360
rect 0 23218 400 23248
rect 3366 23218 3372 23220
rect 0 23158 3372 23218
rect 0 23128 400 23158
rect 3366 23156 3372 23158
rect 3436 23156 3442 23220
rect 2846 22880 3162 22881
rect 2846 22816 2852 22880
rect 2916 22816 2932 22880
rect 2996 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3162 22880
rect 2846 22815 3162 22816
rect 5846 22880 6162 22881
rect 5846 22816 5852 22880
rect 5916 22816 5932 22880
rect 5996 22816 6012 22880
rect 6076 22816 6092 22880
rect 6156 22816 6162 22880
rect 5846 22815 6162 22816
rect 8846 22880 9162 22881
rect 8846 22816 8852 22880
rect 8916 22816 8932 22880
rect 8996 22816 9012 22880
rect 9076 22816 9092 22880
rect 9156 22816 9162 22880
rect 8846 22815 9162 22816
rect 11846 22880 12162 22881
rect 11846 22816 11852 22880
rect 11916 22816 11932 22880
rect 11996 22816 12012 22880
rect 12076 22816 12092 22880
rect 12156 22816 12162 22880
rect 11846 22815 12162 22816
rect 14846 22880 15162 22881
rect 14846 22816 14852 22880
rect 14916 22816 14932 22880
rect 14996 22816 15012 22880
rect 15076 22816 15092 22880
rect 15156 22816 15162 22880
rect 14846 22815 15162 22816
rect 17846 22880 18162 22881
rect 17846 22816 17852 22880
rect 17916 22816 17932 22880
rect 17996 22816 18012 22880
rect 18076 22816 18092 22880
rect 18156 22816 18162 22880
rect 17846 22815 18162 22816
rect 20846 22880 21162 22881
rect 20846 22816 20852 22880
rect 20916 22816 20932 22880
rect 20996 22816 21012 22880
rect 21076 22816 21092 22880
rect 21156 22816 21162 22880
rect 20846 22815 21162 22816
rect 23846 22880 24162 22881
rect 23846 22816 23852 22880
rect 23916 22816 23932 22880
rect 23996 22816 24012 22880
rect 24076 22816 24092 22880
rect 24156 22816 24162 22880
rect 23846 22815 24162 22816
rect 1346 22336 1662 22337
rect 1346 22272 1352 22336
rect 1416 22272 1432 22336
rect 1496 22272 1512 22336
rect 1576 22272 1592 22336
rect 1656 22272 1662 22336
rect 1346 22271 1662 22272
rect 4346 22336 4662 22337
rect 4346 22272 4352 22336
rect 4416 22272 4432 22336
rect 4496 22272 4512 22336
rect 4576 22272 4592 22336
rect 4656 22272 4662 22336
rect 4346 22271 4662 22272
rect 7346 22336 7662 22337
rect 7346 22272 7352 22336
rect 7416 22272 7432 22336
rect 7496 22272 7512 22336
rect 7576 22272 7592 22336
rect 7656 22272 7662 22336
rect 7346 22271 7662 22272
rect 10346 22336 10662 22337
rect 10346 22272 10352 22336
rect 10416 22272 10432 22336
rect 10496 22272 10512 22336
rect 10576 22272 10592 22336
rect 10656 22272 10662 22336
rect 10346 22271 10662 22272
rect 13346 22336 13662 22337
rect 13346 22272 13352 22336
rect 13416 22272 13432 22336
rect 13496 22272 13512 22336
rect 13576 22272 13592 22336
rect 13656 22272 13662 22336
rect 13346 22271 13662 22272
rect 16346 22336 16662 22337
rect 16346 22272 16352 22336
rect 16416 22272 16432 22336
rect 16496 22272 16512 22336
rect 16576 22272 16592 22336
rect 16656 22272 16662 22336
rect 16346 22271 16662 22272
rect 19346 22336 19662 22337
rect 19346 22272 19352 22336
rect 19416 22272 19432 22336
rect 19496 22272 19512 22336
rect 19576 22272 19592 22336
rect 19656 22272 19662 22336
rect 19346 22271 19662 22272
rect 22346 22336 22662 22337
rect 22346 22272 22352 22336
rect 22416 22272 22432 22336
rect 22496 22272 22512 22336
rect 22576 22272 22592 22336
rect 22656 22272 22662 22336
rect 22346 22271 22662 22272
rect 5165 21994 5231 21997
rect 7649 21994 7715 21997
rect 11237 21994 11303 21997
rect 5165 21992 11303 21994
rect 5165 21936 5170 21992
rect 5226 21936 7654 21992
rect 7710 21936 11242 21992
rect 11298 21936 11303 21992
rect 5165 21934 11303 21936
rect 5165 21931 5231 21934
rect 7649 21931 7715 21934
rect 11237 21931 11303 21934
rect 2846 21792 3162 21793
rect 2846 21728 2852 21792
rect 2916 21728 2932 21792
rect 2996 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3162 21792
rect 2846 21727 3162 21728
rect 5846 21792 6162 21793
rect 5846 21728 5852 21792
rect 5916 21728 5932 21792
rect 5996 21728 6012 21792
rect 6076 21728 6092 21792
rect 6156 21728 6162 21792
rect 5846 21727 6162 21728
rect 8846 21792 9162 21793
rect 8846 21728 8852 21792
rect 8916 21728 8932 21792
rect 8996 21728 9012 21792
rect 9076 21728 9092 21792
rect 9156 21728 9162 21792
rect 8846 21727 9162 21728
rect 11846 21792 12162 21793
rect 11846 21728 11852 21792
rect 11916 21728 11932 21792
rect 11996 21728 12012 21792
rect 12076 21728 12092 21792
rect 12156 21728 12162 21792
rect 11846 21727 12162 21728
rect 14846 21792 15162 21793
rect 14846 21728 14852 21792
rect 14916 21728 14932 21792
rect 14996 21728 15012 21792
rect 15076 21728 15092 21792
rect 15156 21728 15162 21792
rect 14846 21727 15162 21728
rect 17846 21792 18162 21793
rect 17846 21728 17852 21792
rect 17916 21728 17932 21792
rect 17996 21728 18012 21792
rect 18076 21728 18092 21792
rect 18156 21728 18162 21792
rect 17846 21727 18162 21728
rect 20846 21792 21162 21793
rect 20846 21728 20852 21792
rect 20916 21728 20932 21792
rect 20996 21728 21012 21792
rect 21076 21728 21092 21792
rect 21156 21728 21162 21792
rect 20846 21727 21162 21728
rect 23846 21792 24162 21793
rect 23846 21728 23852 21792
rect 23916 21728 23932 21792
rect 23996 21728 24012 21792
rect 24076 21728 24092 21792
rect 24156 21728 24162 21792
rect 23846 21727 24162 21728
rect 1346 21248 1662 21249
rect 1346 21184 1352 21248
rect 1416 21184 1432 21248
rect 1496 21184 1512 21248
rect 1576 21184 1592 21248
rect 1656 21184 1662 21248
rect 1346 21183 1662 21184
rect 4346 21248 4662 21249
rect 4346 21184 4352 21248
rect 4416 21184 4432 21248
rect 4496 21184 4512 21248
rect 4576 21184 4592 21248
rect 4656 21184 4662 21248
rect 4346 21183 4662 21184
rect 7346 21248 7662 21249
rect 7346 21184 7352 21248
rect 7416 21184 7432 21248
rect 7496 21184 7512 21248
rect 7576 21184 7592 21248
rect 7656 21184 7662 21248
rect 7346 21183 7662 21184
rect 10346 21248 10662 21249
rect 10346 21184 10352 21248
rect 10416 21184 10432 21248
rect 10496 21184 10512 21248
rect 10576 21184 10592 21248
rect 10656 21184 10662 21248
rect 10346 21183 10662 21184
rect 13346 21248 13662 21249
rect 13346 21184 13352 21248
rect 13416 21184 13432 21248
rect 13496 21184 13512 21248
rect 13576 21184 13592 21248
rect 13656 21184 13662 21248
rect 13346 21183 13662 21184
rect 16346 21248 16662 21249
rect 16346 21184 16352 21248
rect 16416 21184 16432 21248
rect 16496 21184 16512 21248
rect 16576 21184 16592 21248
rect 16656 21184 16662 21248
rect 16346 21183 16662 21184
rect 19346 21248 19662 21249
rect 19346 21184 19352 21248
rect 19416 21184 19432 21248
rect 19496 21184 19512 21248
rect 19576 21184 19592 21248
rect 19656 21184 19662 21248
rect 19346 21183 19662 21184
rect 22346 21248 22662 21249
rect 22346 21184 22352 21248
rect 22416 21184 22432 21248
rect 22496 21184 22512 21248
rect 22576 21184 22592 21248
rect 22656 21184 22662 21248
rect 22346 21183 22662 21184
rect 23565 21178 23631 21181
rect 24780 21178 25180 21208
rect 23565 21176 25180 21178
rect 23565 21120 23570 21176
rect 23626 21120 25180 21176
rect 23565 21118 25180 21120
rect 23565 21115 23631 21118
rect 24780 21088 25180 21118
rect 13629 21042 13695 21045
rect 15101 21042 15167 21045
rect 13629 21040 15167 21042
rect 13629 20984 13634 21040
rect 13690 20984 15106 21040
rect 15162 20984 15167 21040
rect 13629 20982 15167 20984
rect 13629 20979 13695 20982
rect 15101 20979 15167 20982
rect 2846 20704 3162 20705
rect 2846 20640 2852 20704
rect 2916 20640 2932 20704
rect 2996 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3162 20704
rect 2846 20639 3162 20640
rect 5846 20704 6162 20705
rect 5846 20640 5852 20704
rect 5916 20640 5932 20704
rect 5996 20640 6012 20704
rect 6076 20640 6092 20704
rect 6156 20640 6162 20704
rect 5846 20639 6162 20640
rect 8846 20704 9162 20705
rect 8846 20640 8852 20704
rect 8916 20640 8932 20704
rect 8996 20640 9012 20704
rect 9076 20640 9092 20704
rect 9156 20640 9162 20704
rect 8846 20639 9162 20640
rect 11846 20704 12162 20705
rect 11846 20640 11852 20704
rect 11916 20640 11932 20704
rect 11996 20640 12012 20704
rect 12076 20640 12092 20704
rect 12156 20640 12162 20704
rect 11846 20639 12162 20640
rect 14846 20704 15162 20705
rect 14846 20640 14852 20704
rect 14916 20640 14932 20704
rect 14996 20640 15012 20704
rect 15076 20640 15092 20704
rect 15156 20640 15162 20704
rect 14846 20639 15162 20640
rect 17846 20704 18162 20705
rect 17846 20640 17852 20704
rect 17916 20640 17932 20704
rect 17996 20640 18012 20704
rect 18076 20640 18092 20704
rect 18156 20640 18162 20704
rect 17846 20639 18162 20640
rect 20846 20704 21162 20705
rect 20846 20640 20852 20704
rect 20916 20640 20932 20704
rect 20996 20640 21012 20704
rect 21076 20640 21092 20704
rect 21156 20640 21162 20704
rect 20846 20639 21162 20640
rect 23846 20704 24162 20705
rect 23846 20640 23852 20704
rect 23916 20640 23932 20704
rect 23996 20640 24012 20704
rect 24076 20640 24092 20704
rect 24156 20640 24162 20704
rect 23846 20639 24162 20640
rect 1346 20160 1662 20161
rect 1346 20096 1352 20160
rect 1416 20096 1432 20160
rect 1496 20096 1512 20160
rect 1576 20096 1592 20160
rect 1656 20096 1662 20160
rect 1346 20095 1662 20096
rect 4346 20160 4662 20161
rect 4346 20096 4352 20160
rect 4416 20096 4432 20160
rect 4496 20096 4512 20160
rect 4576 20096 4592 20160
rect 4656 20096 4662 20160
rect 4346 20095 4662 20096
rect 7346 20160 7662 20161
rect 7346 20096 7352 20160
rect 7416 20096 7432 20160
rect 7496 20096 7512 20160
rect 7576 20096 7592 20160
rect 7656 20096 7662 20160
rect 7346 20095 7662 20096
rect 10346 20160 10662 20161
rect 10346 20096 10352 20160
rect 10416 20096 10432 20160
rect 10496 20096 10512 20160
rect 10576 20096 10592 20160
rect 10656 20096 10662 20160
rect 10346 20095 10662 20096
rect 13346 20160 13662 20161
rect 13346 20096 13352 20160
rect 13416 20096 13432 20160
rect 13496 20096 13512 20160
rect 13576 20096 13592 20160
rect 13656 20096 13662 20160
rect 13346 20095 13662 20096
rect 16346 20160 16662 20161
rect 16346 20096 16352 20160
rect 16416 20096 16432 20160
rect 16496 20096 16512 20160
rect 16576 20096 16592 20160
rect 16656 20096 16662 20160
rect 16346 20095 16662 20096
rect 19346 20160 19662 20161
rect 19346 20096 19352 20160
rect 19416 20096 19432 20160
rect 19496 20096 19512 20160
rect 19576 20096 19592 20160
rect 19656 20096 19662 20160
rect 19346 20095 19662 20096
rect 22346 20160 22662 20161
rect 22346 20096 22352 20160
rect 22416 20096 22432 20160
rect 22496 20096 22512 20160
rect 22576 20096 22592 20160
rect 22656 20096 22662 20160
rect 22346 20095 22662 20096
rect 23657 19818 23723 19821
rect 24780 19818 25180 19848
rect 23657 19816 25180 19818
rect 23657 19760 23662 19816
rect 23718 19760 25180 19816
rect 23657 19758 25180 19760
rect 23657 19755 23723 19758
rect 24780 19728 25180 19758
rect 2846 19616 3162 19617
rect 2846 19552 2852 19616
rect 2916 19552 2932 19616
rect 2996 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3162 19616
rect 2846 19551 3162 19552
rect 5846 19616 6162 19617
rect 5846 19552 5852 19616
rect 5916 19552 5932 19616
rect 5996 19552 6012 19616
rect 6076 19552 6092 19616
rect 6156 19552 6162 19616
rect 5846 19551 6162 19552
rect 8846 19616 9162 19617
rect 8846 19552 8852 19616
rect 8916 19552 8932 19616
rect 8996 19552 9012 19616
rect 9076 19552 9092 19616
rect 9156 19552 9162 19616
rect 8846 19551 9162 19552
rect 11846 19616 12162 19617
rect 11846 19552 11852 19616
rect 11916 19552 11932 19616
rect 11996 19552 12012 19616
rect 12076 19552 12092 19616
rect 12156 19552 12162 19616
rect 11846 19551 12162 19552
rect 14846 19616 15162 19617
rect 14846 19552 14852 19616
rect 14916 19552 14932 19616
rect 14996 19552 15012 19616
rect 15076 19552 15092 19616
rect 15156 19552 15162 19616
rect 14846 19551 15162 19552
rect 17846 19616 18162 19617
rect 17846 19552 17852 19616
rect 17916 19552 17932 19616
rect 17996 19552 18012 19616
rect 18076 19552 18092 19616
rect 18156 19552 18162 19616
rect 17846 19551 18162 19552
rect 20846 19616 21162 19617
rect 20846 19552 20852 19616
rect 20916 19552 20932 19616
rect 20996 19552 21012 19616
rect 21076 19552 21092 19616
rect 21156 19552 21162 19616
rect 20846 19551 21162 19552
rect 23846 19616 24162 19617
rect 23846 19552 23852 19616
rect 23916 19552 23932 19616
rect 23996 19552 24012 19616
rect 24076 19552 24092 19616
rect 24156 19552 24162 19616
rect 23846 19551 24162 19552
rect 0 19138 400 19168
rect 1209 19138 1275 19141
rect 0 19136 1275 19138
rect 0 19080 1214 19136
rect 1270 19080 1275 19136
rect 0 19078 1275 19080
rect 0 19048 400 19078
rect 1209 19075 1275 19078
rect 23565 19138 23631 19141
rect 24780 19138 25180 19168
rect 23565 19136 25180 19138
rect 23565 19080 23570 19136
rect 23626 19080 25180 19136
rect 23565 19078 25180 19080
rect 23565 19075 23631 19078
rect 1346 19072 1662 19073
rect 1346 19008 1352 19072
rect 1416 19008 1432 19072
rect 1496 19008 1512 19072
rect 1576 19008 1592 19072
rect 1656 19008 1662 19072
rect 1346 19007 1662 19008
rect 4346 19072 4662 19073
rect 4346 19008 4352 19072
rect 4416 19008 4432 19072
rect 4496 19008 4512 19072
rect 4576 19008 4592 19072
rect 4656 19008 4662 19072
rect 4346 19007 4662 19008
rect 7346 19072 7662 19073
rect 7346 19008 7352 19072
rect 7416 19008 7432 19072
rect 7496 19008 7512 19072
rect 7576 19008 7592 19072
rect 7656 19008 7662 19072
rect 7346 19007 7662 19008
rect 10346 19072 10662 19073
rect 10346 19008 10352 19072
rect 10416 19008 10432 19072
rect 10496 19008 10512 19072
rect 10576 19008 10592 19072
rect 10656 19008 10662 19072
rect 10346 19007 10662 19008
rect 13346 19072 13662 19073
rect 13346 19008 13352 19072
rect 13416 19008 13432 19072
rect 13496 19008 13512 19072
rect 13576 19008 13592 19072
rect 13656 19008 13662 19072
rect 13346 19007 13662 19008
rect 16346 19072 16662 19073
rect 16346 19008 16352 19072
rect 16416 19008 16432 19072
rect 16496 19008 16512 19072
rect 16576 19008 16592 19072
rect 16656 19008 16662 19072
rect 16346 19007 16662 19008
rect 19346 19072 19662 19073
rect 19346 19008 19352 19072
rect 19416 19008 19432 19072
rect 19496 19008 19512 19072
rect 19576 19008 19592 19072
rect 19656 19008 19662 19072
rect 19346 19007 19662 19008
rect 22346 19072 22662 19073
rect 22346 19008 22352 19072
rect 22416 19008 22432 19072
rect 22496 19008 22512 19072
rect 22576 19008 22592 19072
rect 22656 19008 22662 19072
rect 24780 19048 25180 19078
rect 22346 19007 22662 19008
rect 2846 18528 3162 18529
rect 0 18461 400 18488
rect 2846 18464 2852 18528
rect 2916 18464 2932 18528
rect 2996 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3162 18528
rect 2846 18463 3162 18464
rect 5846 18528 6162 18529
rect 5846 18464 5852 18528
rect 5916 18464 5932 18528
rect 5996 18464 6012 18528
rect 6076 18464 6092 18528
rect 6156 18464 6162 18528
rect 5846 18463 6162 18464
rect 8846 18528 9162 18529
rect 8846 18464 8852 18528
rect 8916 18464 8932 18528
rect 8996 18464 9012 18528
rect 9076 18464 9092 18528
rect 9156 18464 9162 18528
rect 8846 18463 9162 18464
rect 11846 18528 12162 18529
rect 11846 18464 11852 18528
rect 11916 18464 11932 18528
rect 11996 18464 12012 18528
rect 12076 18464 12092 18528
rect 12156 18464 12162 18528
rect 11846 18463 12162 18464
rect 14846 18528 15162 18529
rect 14846 18464 14852 18528
rect 14916 18464 14932 18528
rect 14996 18464 15012 18528
rect 15076 18464 15092 18528
rect 15156 18464 15162 18528
rect 14846 18463 15162 18464
rect 17846 18528 18162 18529
rect 17846 18464 17852 18528
rect 17916 18464 17932 18528
rect 17996 18464 18012 18528
rect 18076 18464 18092 18528
rect 18156 18464 18162 18528
rect 17846 18463 18162 18464
rect 20846 18528 21162 18529
rect 20846 18464 20852 18528
rect 20916 18464 20932 18528
rect 20996 18464 21012 18528
rect 21076 18464 21092 18528
rect 21156 18464 21162 18528
rect 20846 18463 21162 18464
rect 23846 18528 24162 18529
rect 23846 18464 23852 18528
rect 23916 18464 23932 18528
rect 23996 18464 24012 18528
rect 24076 18464 24092 18528
rect 24156 18464 24162 18528
rect 23846 18463 24162 18464
rect 0 18456 447 18461
rect 0 18400 386 18456
rect 442 18400 447 18456
rect 0 18395 447 18400
rect 24301 18458 24367 18461
rect 24780 18458 25180 18488
rect 24301 18456 25180 18458
rect 24301 18400 24306 18456
rect 24362 18400 25180 18456
rect 24301 18398 25180 18400
rect 24301 18395 24367 18398
rect 0 18368 400 18395
rect 24780 18368 25180 18398
rect 10961 18322 11027 18325
rect 13118 18322 13124 18324
rect 10961 18320 13124 18322
rect 10961 18264 10966 18320
rect 11022 18264 13124 18320
rect 10961 18262 13124 18264
rect 10961 18259 11027 18262
rect 13118 18260 13124 18262
rect 13188 18322 13194 18324
rect 16665 18322 16731 18325
rect 13188 18320 20730 18322
rect 13188 18264 16670 18320
rect 16726 18264 20730 18320
rect 13188 18262 20730 18264
rect 13188 18260 13194 18262
rect 16665 18259 16731 18262
rect 1346 17984 1662 17985
rect 1346 17920 1352 17984
rect 1416 17920 1432 17984
rect 1496 17920 1512 17984
rect 1576 17920 1592 17984
rect 1656 17920 1662 17984
rect 1346 17919 1662 17920
rect 4346 17984 4662 17985
rect 4346 17920 4352 17984
rect 4416 17920 4432 17984
rect 4496 17920 4512 17984
rect 4576 17920 4592 17984
rect 4656 17920 4662 17984
rect 4346 17919 4662 17920
rect 7346 17984 7662 17985
rect 7346 17920 7352 17984
rect 7416 17920 7432 17984
rect 7496 17920 7512 17984
rect 7576 17920 7592 17984
rect 7656 17920 7662 17984
rect 7346 17919 7662 17920
rect 10346 17984 10662 17985
rect 10346 17920 10352 17984
rect 10416 17920 10432 17984
rect 10496 17920 10512 17984
rect 10576 17920 10592 17984
rect 10656 17920 10662 17984
rect 10346 17919 10662 17920
rect 13346 17984 13662 17985
rect 13346 17920 13352 17984
rect 13416 17920 13432 17984
rect 13496 17920 13512 17984
rect 13576 17920 13592 17984
rect 13656 17920 13662 17984
rect 13346 17919 13662 17920
rect 16346 17984 16662 17985
rect 16346 17920 16352 17984
rect 16416 17920 16432 17984
rect 16496 17920 16512 17984
rect 16576 17920 16592 17984
rect 16656 17920 16662 17984
rect 16346 17919 16662 17920
rect 19346 17984 19662 17985
rect 19346 17920 19352 17984
rect 19416 17920 19432 17984
rect 19496 17920 19512 17984
rect 19576 17920 19592 17984
rect 19656 17920 19662 17984
rect 19346 17919 19662 17920
rect 20670 17917 20730 18262
rect 22134 18124 22140 18188
rect 22204 18186 22210 18188
rect 22369 18186 22435 18189
rect 22204 18184 22435 18186
rect 22204 18128 22374 18184
rect 22430 18128 22435 18184
rect 22204 18126 22435 18128
rect 22204 18124 22210 18126
rect 22369 18123 22435 18126
rect 22346 17984 22662 17985
rect 22346 17920 22352 17984
rect 22416 17920 22432 17984
rect 22496 17920 22512 17984
rect 22576 17920 22592 17984
rect 22656 17920 22662 17984
rect 22346 17919 22662 17920
rect 20670 17912 20779 17917
rect 20670 17856 20718 17912
rect 20774 17856 20779 17912
rect 20670 17854 20779 17856
rect 20713 17851 20779 17854
rect 23289 17778 23355 17781
rect 24780 17778 25180 17808
rect 23289 17776 25180 17778
rect 23289 17720 23294 17776
rect 23350 17720 25180 17776
rect 23289 17718 25180 17720
rect 23289 17715 23355 17718
rect 24780 17688 25180 17718
rect 14273 17642 14339 17645
rect 14549 17642 14615 17645
rect 14917 17642 14983 17645
rect 14273 17640 14983 17642
rect 14273 17584 14278 17640
rect 14334 17584 14554 17640
rect 14610 17584 14922 17640
rect 14978 17584 14983 17640
rect 14273 17582 14983 17584
rect 14273 17579 14339 17582
rect 14549 17579 14615 17582
rect 14917 17579 14983 17582
rect 2846 17440 3162 17441
rect 2846 17376 2852 17440
rect 2916 17376 2932 17440
rect 2996 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3162 17440
rect 2846 17375 3162 17376
rect 5846 17440 6162 17441
rect 5846 17376 5852 17440
rect 5916 17376 5932 17440
rect 5996 17376 6012 17440
rect 6076 17376 6092 17440
rect 6156 17376 6162 17440
rect 5846 17375 6162 17376
rect 8846 17440 9162 17441
rect 8846 17376 8852 17440
rect 8916 17376 8932 17440
rect 8996 17376 9012 17440
rect 9076 17376 9092 17440
rect 9156 17376 9162 17440
rect 8846 17375 9162 17376
rect 11846 17440 12162 17441
rect 11846 17376 11852 17440
rect 11916 17376 11932 17440
rect 11996 17376 12012 17440
rect 12076 17376 12092 17440
rect 12156 17376 12162 17440
rect 11846 17375 12162 17376
rect 14846 17440 15162 17441
rect 14846 17376 14852 17440
rect 14916 17376 14932 17440
rect 14996 17376 15012 17440
rect 15076 17376 15092 17440
rect 15156 17376 15162 17440
rect 14846 17375 15162 17376
rect 17846 17440 18162 17441
rect 17846 17376 17852 17440
rect 17916 17376 17932 17440
rect 17996 17376 18012 17440
rect 18076 17376 18092 17440
rect 18156 17376 18162 17440
rect 17846 17375 18162 17376
rect 20846 17440 21162 17441
rect 20846 17376 20852 17440
rect 20916 17376 20932 17440
rect 20996 17376 21012 17440
rect 21076 17376 21092 17440
rect 21156 17376 21162 17440
rect 20846 17375 21162 17376
rect 23846 17440 24162 17441
rect 23846 17376 23852 17440
rect 23916 17376 23932 17440
rect 23996 17376 24012 17440
rect 24076 17376 24092 17440
rect 24156 17376 24162 17440
rect 23846 17375 24162 17376
rect 23749 17098 23815 17101
rect 24780 17098 25180 17128
rect 23749 17096 25180 17098
rect 23749 17040 23754 17096
rect 23810 17040 25180 17096
rect 23749 17038 25180 17040
rect 23749 17035 23815 17038
rect 24780 17008 25180 17038
rect 1346 16896 1662 16897
rect 1346 16832 1352 16896
rect 1416 16832 1432 16896
rect 1496 16832 1512 16896
rect 1576 16832 1592 16896
rect 1656 16832 1662 16896
rect 1346 16831 1662 16832
rect 4346 16896 4662 16897
rect 4346 16832 4352 16896
rect 4416 16832 4432 16896
rect 4496 16832 4512 16896
rect 4576 16832 4592 16896
rect 4656 16832 4662 16896
rect 4346 16831 4662 16832
rect 7346 16896 7662 16897
rect 7346 16832 7352 16896
rect 7416 16832 7432 16896
rect 7496 16832 7512 16896
rect 7576 16832 7592 16896
rect 7656 16832 7662 16896
rect 7346 16831 7662 16832
rect 10346 16896 10662 16897
rect 10346 16832 10352 16896
rect 10416 16832 10432 16896
rect 10496 16832 10512 16896
rect 10576 16832 10592 16896
rect 10656 16832 10662 16896
rect 10346 16831 10662 16832
rect 13346 16896 13662 16897
rect 13346 16832 13352 16896
rect 13416 16832 13432 16896
rect 13496 16832 13512 16896
rect 13576 16832 13592 16896
rect 13656 16832 13662 16896
rect 13346 16831 13662 16832
rect 16346 16896 16662 16897
rect 16346 16832 16352 16896
rect 16416 16832 16432 16896
rect 16496 16832 16512 16896
rect 16576 16832 16592 16896
rect 16656 16832 16662 16896
rect 16346 16831 16662 16832
rect 19346 16896 19662 16897
rect 19346 16832 19352 16896
rect 19416 16832 19432 16896
rect 19496 16832 19512 16896
rect 19576 16832 19592 16896
rect 19656 16832 19662 16896
rect 19346 16831 19662 16832
rect 22346 16896 22662 16897
rect 22346 16832 22352 16896
rect 22416 16832 22432 16896
rect 22496 16832 22512 16896
rect 22576 16832 22592 16896
rect 22656 16832 22662 16896
rect 22346 16831 22662 16832
rect 23381 16554 23447 16557
rect 23381 16552 24410 16554
rect 23381 16496 23386 16552
rect 23442 16496 24410 16552
rect 23381 16494 24410 16496
rect 23381 16491 23447 16494
rect 0 16418 400 16448
rect 1301 16418 1367 16421
rect 0 16416 1367 16418
rect 0 16360 1306 16416
rect 1362 16360 1367 16416
rect 0 16358 1367 16360
rect 24350 16418 24410 16494
rect 24780 16418 25180 16448
rect 24350 16358 25180 16418
rect 0 16328 400 16358
rect 1301 16355 1367 16358
rect 2846 16352 3162 16353
rect 2846 16288 2852 16352
rect 2916 16288 2932 16352
rect 2996 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3162 16352
rect 2846 16287 3162 16288
rect 5846 16352 6162 16353
rect 5846 16288 5852 16352
rect 5916 16288 5932 16352
rect 5996 16288 6012 16352
rect 6076 16288 6092 16352
rect 6156 16288 6162 16352
rect 5846 16287 6162 16288
rect 8846 16352 9162 16353
rect 8846 16288 8852 16352
rect 8916 16288 8932 16352
rect 8996 16288 9012 16352
rect 9076 16288 9092 16352
rect 9156 16288 9162 16352
rect 8846 16287 9162 16288
rect 11846 16352 12162 16353
rect 11846 16288 11852 16352
rect 11916 16288 11932 16352
rect 11996 16288 12012 16352
rect 12076 16288 12092 16352
rect 12156 16288 12162 16352
rect 11846 16287 12162 16288
rect 14846 16352 15162 16353
rect 14846 16288 14852 16352
rect 14916 16288 14932 16352
rect 14996 16288 15012 16352
rect 15076 16288 15092 16352
rect 15156 16288 15162 16352
rect 14846 16287 15162 16288
rect 17846 16352 18162 16353
rect 17846 16288 17852 16352
rect 17916 16288 17932 16352
rect 17996 16288 18012 16352
rect 18076 16288 18092 16352
rect 18156 16288 18162 16352
rect 17846 16287 18162 16288
rect 20846 16352 21162 16353
rect 20846 16288 20852 16352
rect 20916 16288 20932 16352
rect 20996 16288 21012 16352
rect 21076 16288 21092 16352
rect 21156 16288 21162 16352
rect 20846 16287 21162 16288
rect 23846 16352 24162 16353
rect 23846 16288 23852 16352
rect 23916 16288 23932 16352
rect 23996 16288 24012 16352
rect 24076 16288 24092 16352
rect 24156 16288 24162 16352
rect 24780 16328 25180 16358
rect 23846 16287 24162 16288
rect 1346 15808 1662 15809
rect 0 15738 400 15768
rect 1346 15744 1352 15808
rect 1416 15744 1432 15808
rect 1496 15744 1512 15808
rect 1576 15744 1592 15808
rect 1656 15744 1662 15808
rect 1346 15743 1662 15744
rect 4346 15808 4662 15809
rect 4346 15744 4352 15808
rect 4416 15744 4432 15808
rect 4496 15744 4512 15808
rect 4576 15744 4592 15808
rect 4656 15744 4662 15808
rect 4346 15743 4662 15744
rect 7346 15808 7662 15809
rect 7346 15744 7352 15808
rect 7416 15744 7432 15808
rect 7496 15744 7512 15808
rect 7576 15744 7592 15808
rect 7656 15744 7662 15808
rect 7346 15743 7662 15744
rect 10346 15808 10662 15809
rect 10346 15744 10352 15808
rect 10416 15744 10432 15808
rect 10496 15744 10512 15808
rect 10576 15744 10592 15808
rect 10656 15744 10662 15808
rect 10346 15743 10662 15744
rect 13346 15808 13662 15809
rect 13346 15744 13352 15808
rect 13416 15744 13432 15808
rect 13496 15744 13512 15808
rect 13576 15744 13592 15808
rect 13656 15744 13662 15808
rect 13346 15743 13662 15744
rect 16346 15808 16662 15809
rect 16346 15744 16352 15808
rect 16416 15744 16432 15808
rect 16496 15744 16512 15808
rect 16576 15744 16592 15808
rect 16656 15744 16662 15808
rect 16346 15743 16662 15744
rect 19346 15808 19662 15809
rect 19346 15744 19352 15808
rect 19416 15744 19432 15808
rect 19496 15744 19512 15808
rect 19576 15744 19592 15808
rect 19656 15744 19662 15808
rect 19346 15743 19662 15744
rect 22346 15808 22662 15809
rect 22346 15744 22352 15808
rect 22416 15744 22432 15808
rect 22496 15744 22512 15808
rect 22576 15744 22592 15808
rect 22656 15744 22662 15808
rect 22346 15743 22662 15744
rect 749 15738 815 15741
rect 0 15736 815 15738
rect 0 15680 754 15736
rect 810 15680 815 15736
rect 0 15678 815 15680
rect 0 15648 400 15678
rect 749 15675 815 15678
rect 23381 15738 23447 15741
rect 24780 15738 25180 15768
rect 23381 15736 25180 15738
rect 23381 15680 23386 15736
rect 23442 15680 25180 15736
rect 23381 15678 25180 15680
rect 23381 15675 23447 15678
rect 24780 15648 25180 15678
rect 19241 15602 19307 15605
rect 22277 15602 22343 15605
rect 19241 15600 22343 15602
rect 19241 15544 19246 15600
rect 19302 15544 22282 15600
rect 22338 15544 22343 15600
rect 19241 15542 22343 15544
rect 19241 15539 19307 15542
rect 22277 15539 22343 15542
rect 2846 15264 3162 15265
rect 2846 15200 2852 15264
rect 2916 15200 2932 15264
rect 2996 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3162 15264
rect 2846 15199 3162 15200
rect 5846 15264 6162 15265
rect 5846 15200 5852 15264
rect 5916 15200 5932 15264
rect 5996 15200 6012 15264
rect 6076 15200 6092 15264
rect 6156 15200 6162 15264
rect 5846 15199 6162 15200
rect 8846 15264 9162 15265
rect 8846 15200 8852 15264
rect 8916 15200 8932 15264
rect 8996 15200 9012 15264
rect 9076 15200 9092 15264
rect 9156 15200 9162 15264
rect 8846 15199 9162 15200
rect 11846 15264 12162 15265
rect 11846 15200 11852 15264
rect 11916 15200 11932 15264
rect 11996 15200 12012 15264
rect 12076 15200 12092 15264
rect 12156 15200 12162 15264
rect 11846 15199 12162 15200
rect 14846 15264 15162 15265
rect 14846 15200 14852 15264
rect 14916 15200 14932 15264
rect 14996 15200 15012 15264
rect 15076 15200 15092 15264
rect 15156 15200 15162 15264
rect 14846 15199 15162 15200
rect 17846 15264 18162 15265
rect 17846 15200 17852 15264
rect 17916 15200 17932 15264
rect 17996 15200 18012 15264
rect 18076 15200 18092 15264
rect 18156 15200 18162 15264
rect 17846 15199 18162 15200
rect 20846 15264 21162 15265
rect 20846 15200 20852 15264
rect 20916 15200 20932 15264
rect 20996 15200 21012 15264
rect 21076 15200 21092 15264
rect 21156 15200 21162 15264
rect 20846 15199 21162 15200
rect 23846 15264 24162 15265
rect 23846 15200 23852 15264
rect 23916 15200 23932 15264
rect 23996 15200 24012 15264
rect 24076 15200 24092 15264
rect 24156 15200 24162 15264
rect 23846 15199 24162 15200
rect 0 15058 400 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 400 14998
rect 1393 14995 1459 14998
rect 21541 15058 21607 15061
rect 24780 15058 25180 15088
rect 21541 15056 25180 15058
rect 21541 15000 21546 15056
rect 21602 15000 25180 15056
rect 21541 14998 25180 15000
rect 21541 14995 21607 14998
rect 24780 14968 25180 14998
rect 1346 14720 1662 14721
rect 1346 14656 1352 14720
rect 1416 14656 1432 14720
rect 1496 14656 1512 14720
rect 1576 14656 1592 14720
rect 1656 14656 1662 14720
rect 1346 14655 1662 14656
rect 4346 14720 4662 14721
rect 4346 14656 4352 14720
rect 4416 14656 4432 14720
rect 4496 14656 4512 14720
rect 4576 14656 4592 14720
rect 4656 14656 4662 14720
rect 4346 14655 4662 14656
rect 7346 14720 7662 14721
rect 7346 14656 7352 14720
rect 7416 14656 7432 14720
rect 7496 14656 7512 14720
rect 7576 14656 7592 14720
rect 7656 14656 7662 14720
rect 7346 14655 7662 14656
rect 10346 14720 10662 14721
rect 10346 14656 10352 14720
rect 10416 14656 10432 14720
rect 10496 14656 10512 14720
rect 10576 14656 10592 14720
rect 10656 14656 10662 14720
rect 10346 14655 10662 14656
rect 13346 14720 13662 14721
rect 13346 14656 13352 14720
rect 13416 14656 13432 14720
rect 13496 14656 13512 14720
rect 13576 14656 13592 14720
rect 13656 14656 13662 14720
rect 13346 14655 13662 14656
rect 16346 14720 16662 14721
rect 16346 14656 16352 14720
rect 16416 14656 16432 14720
rect 16496 14656 16512 14720
rect 16576 14656 16592 14720
rect 16656 14656 16662 14720
rect 16346 14655 16662 14656
rect 19346 14720 19662 14721
rect 19346 14656 19352 14720
rect 19416 14656 19432 14720
rect 19496 14656 19512 14720
rect 19576 14656 19592 14720
rect 19656 14656 19662 14720
rect 19346 14655 19662 14656
rect 22346 14720 22662 14721
rect 22346 14656 22352 14720
rect 22416 14656 22432 14720
rect 22496 14656 22512 14720
rect 22576 14656 22592 14720
rect 22656 14656 22662 14720
rect 22346 14655 22662 14656
rect 0 14378 400 14408
rect 749 14378 815 14381
rect 0 14376 815 14378
rect 0 14320 754 14376
rect 810 14320 815 14376
rect 0 14318 815 14320
rect 0 14288 400 14318
rect 749 14315 815 14318
rect 23565 14378 23631 14381
rect 24780 14378 25180 14408
rect 23565 14376 25180 14378
rect 23565 14320 23570 14376
rect 23626 14320 25180 14376
rect 23565 14318 25180 14320
rect 23565 14315 23631 14318
rect 24780 14288 25180 14318
rect 2846 14176 3162 14177
rect 2846 14112 2852 14176
rect 2916 14112 2932 14176
rect 2996 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3162 14176
rect 2846 14111 3162 14112
rect 5846 14176 6162 14177
rect 5846 14112 5852 14176
rect 5916 14112 5932 14176
rect 5996 14112 6012 14176
rect 6076 14112 6092 14176
rect 6156 14112 6162 14176
rect 5846 14111 6162 14112
rect 8846 14176 9162 14177
rect 8846 14112 8852 14176
rect 8916 14112 8932 14176
rect 8996 14112 9012 14176
rect 9076 14112 9092 14176
rect 9156 14112 9162 14176
rect 8846 14111 9162 14112
rect 11846 14176 12162 14177
rect 11846 14112 11852 14176
rect 11916 14112 11932 14176
rect 11996 14112 12012 14176
rect 12076 14112 12092 14176
rect 12156 14112 12162 14176
rect 11846 14111 12162 14112
rect 14846 14176 15162 14177
rect 14846 14112 14852 14176
rect 14916 14112 14932 14176
rect 14996 14112 15012 14176
rect 15076 14112 15092 14176
rect 15156 14112 15162 14176
rect 14846 14111 15162 14112
rect 17846 14176 18162 14177
rect 17846 14112 17852 14176
rect 17916 14112 17932 14176
rect 17996 14112 18012 14176
rect 18076 14112 18092 14176
rect 18156 14112 18162 14176
rect 17846 14111 18162 14112
rect 20846 14176 21162 14177
rect 20846 14112 20852 14176
rect 20916 14112 20932 14176
rect 20996 14112 21012 14176
rect 21076 14112 21092 14176
rect 21156 14112 21162 14176
rect 20846 14111 21162 14112
rect 23846 14176 24162 14177
rect 23846 14112 23852 14176
rect 23916 14112 23932 14176
rect 23996 14112 24012 14176
rect 24076 14112 24092 14176
rect 24156 14112 24162 14176
rect 23846 14111 24162 14112
rect 3366 13908 3372 13972
rect 3436 13970 3442 13972
rect 12525 13970 12591 13973
rect 3436 13968 12591 13970
rect 3436 13912 12530 13968
rect 12586 13912 12591 13968
rect 3436 13910 12591 13912
rect 3436 13908 3442 13910
rect 12525 13907 12591 13910
rect 13118 13908 13124 13972
rect 13188 13970 13194 13972
rect 13721 13970 13787 13973
rect 13188 13968 13787 13970
rect 13188 13912 13726 13968
rect 13782 13912 13787 13968
rect 13188 13910 13787 13912
rect 13188 13908 13194 13910
rect 13721 13907 13787 13910
rect 0 13698 400 13728
rect 1209 13698 1275 13701
rect 0 13696 1275 13698
rect 0 13640 1214 13696
rect 1270 13640 1275 13696
rect 0 13638 1275 13640
rect 0 13608 400 13638
rect 1209 13635 1275 13638
rect 22093 13700 22159 13701
rect 22093 13696 22140 13700
rect 22204 13698 22210 13700
rect 23657 13698 23723 13701
rect 24780 13698 25180 13728
rect 22093 13640 22098 13696
rect 22093 13636 22140 13640
rect 22204 13638 22250 13698
rect 23657 13696 25180 13698
rect 23657 13640 23662 13696
rect 23718 13640 25180 13696
rect 23657 13638 25180 13640
rect 22204 13636 22210 13638
rect 22093 13635 22159 13636
rect 23657 13635 23723 13638
rect 1346 13632 1662 13633
rect 1346 13568 1352 13632
rect 1416 13568 1432 13632
rect 1496 13568 1512 13632
rect 1576 13568 1592 13632
rect 1656 13568 1662 13632
rect 1346 13567 1662 13568
rect 4346 13632 4662 13633
rect 4346 13568 4352 13632
rect 4416 13568 4432 13632
rect 4496 13568 4512 13632
rect 4576 13568 4592 13632
rect 4656 13568 4662 13632
rect 4346 13567 4662 13568
rect 7346 13632 7662 13633
rect 7346 13568 7352 13632
rect 7416 13568 7432 13632
rect 7496 13568 7512 13632
rect 7576 13568 7592 13632
rect 7656 13568 7662 13632
rect 7346 13567 7662 13568
rect 10346 13632 10662 13633
rect 10346 13568 10352 13632
rect 10416 13568 10432 13632
rect 10496 13568 10512 13632
rect 10576 13568 10592 13632
rect 10656 13568 10662 13632
rect 10346 13567 10662 13568
rect 13346 13632 13662 13633
rect 13346 13568 13352 13632
rect 13416 13568 13432 13632
rect 13496 13568 13512 13632
rect 13576 13568 13592 13632
rect 13656 13568 13662 13632
rect 13346 13567 13662 13568
rect 16346 13632 16662 13633
rect 16346 13568 16352 13632
rect 16416 13568 16432 13632
rect 16496 13568 16512 13632
rect 16576 13568 16592 13632
rect 16656 13568 16662 13632
rect 16346 13567 16662 13568
rect 19346 13632 19662 13633
rect 19346 13568 19352 13632
rect 19416 13568 19432 13632
rect 19496 13568 19512 13632
rect 19576 13568 19592 13632
rect 19656 13568 19662 13632
rect 19346 13567 19662 13568
rect 22346 13632 22662 13633
rect 22346 13568 22352 13632
rect 22416 13568 22432 13632
rect 22496 13568 22512 13632
rect 22576 13568 22592 13632
rect 22656 13568 22662 13632
rect 24780 13608 25180 13638
rect 22346 13567 22662 13568
rect 2846 13088 3162 13089
rect 0 13018 400 13048
rect 2846 13024 2852 13088
rect 2916 13024 2932 13088
rect 2996 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3162 13088
rect 2846 13023 3162 13024
rect 5846 13088 6162 13089
rect 5846 13024 5852 13088
rect 5916 13024 5932 13088
rect 5996 13024 6012 13088
rect 6076 13024 6092 13088
rect 6156 13024 6162 13088
rect 5846 13023 6162 13024
rect 8846 13088 9162 13089
rect 8846 13024 8852 13088
rect 8916 13024 8932 13088
rect 8996 13024 9012 13088
rect 9076 13024 9092 13088
rect 9156 13024 9162 13088
rect 8846 13023 9162 13024
rect 11846 13088 12162 13089
rect 11846 13024 11852 13088
rect 11916 13024 11932 13088
rect 11996 13024 12012 13088
rect 12076 13024 12092 13088
rect 12156 13024 12162 13088
rect 11846 13023 12162 13024
rect 14846 13088 15162 13089
rect 14846 13024 14852 13088
rect 14916 13024 14932 13088
rect 14996 13024 15012 13088
rect 15076 13024 15092 13088
rect 15156 13024 15162 13088
rect 14846 13023 15162 13024
rect 17846 13088 18162 13089
rect 17846 13024 17852 13088
rect 17916 13024 17932 13088
rect 17996 13024 18012 13088
rect 18076 13024 18092 13088
rect 18156 13024 18162 13088
rect 17846 13023 18162 13024
rect 20846 13088 21162 13089
rect 20846 13024 20852 13088
rect 20916 13024 20932 13088
rect 20996 13024 21012 13088
rect 21076 13024 21092 13088
rect 21156 13024 21162 13088
rect 20846 13023 21162 13024
rect 23846 13088 24162 13089
rect 23846 13024 23852 13088
rect 23916 13024 23932 13088
rect 23996 13024 24012 13088
rect 24076 13024 24092 13088
rect 24156 13024 24162 13088
rect 23846 13023 24162 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 400 12958
rect 1301 12955 1367 12958
rect 24301 13018 24367 13021
rect 24780 13018 25180 13048
rect 24301 13016 25180 13018
rect 24301 12960 24306 13016
rect 24362 12960 25180 13016
rect 24301 12958 25180 12960
rect 24301 12955 24367 12958
rect 24780 12928 25180 12958
rect 3877 12746 3943 12749
rect 6177 12746 6243 12749
rect 3877 12744 6243 12746
rect 3877 12688 3882 12744
rect 3938 12688 6182 12744
rect 6238 12688 6243 12744
rect 3877 12686 6243 12688
rect 3877 12683 3943 12686
rect 6177 12683 6243 12686
rect 1346 12544 1662 12545
rect 1346 12480 1352 12544
rect 1416 12480 1432 12544
rect 1496 12480 1512 12544
rect 1576 12480 1592 12544
rect 1656 12480 1662 12544
rect 1346 12479 1662 12480
rect 4346 12544 4662 12545
rect 4346 12480 4352 12544
rect 4416 12480 4432 12544
rect 4496 12480 4512 12544
rect 4576 12480 4592 12544
rect 4656 12480 4662 12544
rect 4346 12479 4662 12480
rect 7346 12544 7662 12545
rect 7346 12480 7352 12544
rect 7416 12480 7432 12544
rect 7496 12480 7512 12544
rect 7576 12480 7592 12544
rect 7656 12480 7662 12544
rect 7346 12479 7662 12480
rect 10346 12544 10662 12545
rect 10346 12480 10352 12544
rect 10416 12480 10432 12544
rect 10496 12480 10512 12544
rect 10576 12480 10592 12544
rect 10656 12480 10662 12544
rect 10346 12479 10662 12480
rect 13346 12544 13662 12545
rect 13346 12480 13352 12544
rect 13416 12480 13432 12544
rect 13496 12480 13512 12544
rect 13576 12480 13592 12544
rect 13656 12480 13662 12544
rect 13346 12479 13662 12480
rect 16346 12544 16662 12545
rect 16346 12480 16352 12544
rect 16416 12480 16432 12544
rect 16496 12480 16512 12544
rect 16576 12480 16592 12544
rect 16656 12480 16662 12544
rect 16346 12479 16662 12480
rect 19346 12544 19662 12545
rect 19346 12480 19352 12544
rect 19416 12480 19432 12544
rect 19496 12480 19512 12544
rect 19576 12480 19592 12544
rect 19656 12480 19662 12544
rect 19346 12479 19662 12480
rect 22346 12544 22662 12545
rect 22346 12480 22352 12544
rect 22416 12480 22432 12544
rect 22496 12480 22512 12544
rect 22576 12480 22592 12544
rect 22656 12480 22662 12544
rect 22346 12479 22662 12480
rect 0 12341 400 12368
rect 0 12336 447 12341
rect 0 12280 386 12336
rect 442 12280 447 12336
rect 0 12275 447 12280
rect 23565 12338 23631 12341
rect 24780 12338 25180 12368
rect 23565 12336 25180 12338
rect 23565 12280 23570 12336
rect 23626 12280 25180 12336
rect 23565 12278 25180 12280
rect 23565 12275 23631 12278
rect 0 12248 400 12275
rect 24780 12248 25180 12278
rect 2846 12000 3162 12001
rect 2846 11936 2852 12000
rect 2916 11936 2932 12000
rect 2996 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3162 12000
rect 2846 11935 3162 11936
rect 5846 12000 6162 12001
rect 5846 11936 5852 12000
rect 5916 11936 5932 12000
rect 5996 11936 6012 12000
rect 6076 11936 6092 12000
rect 6156 11936 6162 12000
rect 5846 11935 6162 11936
rect 8846 12000 9162 12001
rect 8846 11936 8852 12000
rect 8916 11936 8932 12000
rect 8996 11936 9012 12000
rect 9076 11936 9092 12000
rect 9156 11936 9162 12000
rect 8846 11935 9162 11936
rect 11846 12000 12162 12001
rect 11846 11936 11852 12000
rect 11916 11936 11932 12000
rect 11996 11936 12012 12000
rect 12076 11936 12092 12000
rect 12156 11936 12162 12000
rect 11846 11935 12162 11936
rect 14846 12000 15162 12001
rect 14846 11936 14852 12000
rect 14916 11936 14932 12000
rect 14996 11936 15012 12000
rect 15076 11936 15092 12000
rect 15156 11936 15162 12000
rect 14846 11935 15162 11936
rect 17846 12000 18162 12001
rect 17846 11936 17852 12000
rect 17916 11936 17932 12000
rect 17996 11936 18012 12000
rect 18076 11936 18092 12000
rect 18156 11936 18162 12000
rect 17846 11935 18162 11936
rect 20846 12000 21162 12001
rect 20846 11936 20852 12000
rect 20916 11936 20932 12000
rect 20996 11936 21012 12000
rect 21076 11936 21092 12000
rect 21156 11936 21162 12000
rect 20846 11935 21162 11936
rect 23846 12000 24162 12001
rect 23846 11936 23852 12000
rect 23916 11936 23932 12000
rect 23996 11936 24012 12000
rect 24076 11936 24092 12000
rect 24156 11936 24162 12000
rect 23846 11935 24162 11936
rect 0 11661 400 11688
rect 0 11656 447 11661
rect 0 11600 386 11656
rect 442 11600 447 11656
rect 0 11595 447 11600
rect 23473 11658 23539 11661
rect 24780 11658 25180 11688
rect 23473 11656 25180 11658
rect 23473 11600 23478 11656
rect 23534 11600 25180 11656
rect 23473 11598 25180 11600
rect 23473 11595 23539 11598
rect 0 11568 400 11595
rect 24780 11568 25180 11598
rect 1346 11456 1662 11457
rect 1346 11392 1352 11456
rect 1416 11392 1432 11456
rect 1496 11392 1512 11456
rect 1576 11392 1592 11456
rect 1656 11392 1662 11456
rect 1346 11391 1662 11392
rect 4346 11456 4662 11457
rect 4346 11392 4352 11456
rect 4416 11392 4432 11456
rect 4496 11392 4512 11456
rect 4576 11392 4592 11456
rect 4656 11392 4662 11456
rect 4346 11391 4662 11392
rect 7346 11456 7662 11457
rect 7346 11392 7352 11456
rect 7416 11392 7432 11456
rect 7496 11392 7512 11456
rect 7576 11392 7592 11456
rect 7656 11392 7662 11456
rect 7346 11391 7662 11392
rect 10346 11456 10662 11457
rect 10346 11392 10352 11456
rect 10416 11392 10432 11456
rect 10496 11392 10512 11456
rect 10576 11392 10592 11456
rect 10656 11392 10662 11456
rect 10346 11391 10662 11392
rect 13346 11456 13662 11457
rect 13346 11392 13352 11456
rect 13416 11392 13432 11456
rect 13496 11392 13512 11456
rect 13576 11392 13592 11456
rect 13656 11392 13662 11456
rect 13346 11391 13662 11392
rect 16346 11456 16662 11457
rect 16346 11392 16352 11456
rect 16416 11392 16432 11456
rect 16496 11392 16512 11456
rect 16576 11392 16592 11456
rect 16656 11392 16662 11456
rect 16346 11391 16662 11392
rect 19346 11456 19662 11457
rect 19346 11392 19352 11456
rect 19416 11392 19432 11456
rect 19496 11392 19512 11456
rect 19576 11392 19592 11456
rect 19656 11392 19662 11456
rect 19346 11391 19662 11392
rect 22346 11456 22662 11457
rect 22346 11392 22352 11456
rect 22416 11392 22432 11456
rect 22496 11392 22512 11456
rect 22576 11392 22592 11456
rect 22656 11392 22662 11456
rect 22346 11391 22662 11392
rect 8937 11114 9003 11117
rect 13118 11114 13124 11116
rect 8937 11112 13124 11114
rect 8937 11056 8942 11112
rect 8998 11056 13124 11112
rect 8937 11054 13124 11056
rect 8937 11051 9003 11054
rect 13118 11052 13124 11054
rect 13188 11114 13194 11116
rect 14365 11114 14431 11117
rect 13188 11112 14431 11114
rect 13188 11056 14370 11112
rect 14426 11056 14431 11112
rect 13188 11054 14431 11056
rect 13188 11052 13194 11054
rect 14365 11051 14431 11054
rect 0 10978 400 11008
rect 1485 10978 1551 10981
rect 24780 10978 25180 11008
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 400 10918
rect 1485 10915 1551 10918
rect 24350 10918 25180 10978
rect 2846 10912 3162 10913
rect 2846 10848 2852 10912
rect 2916 10848 2932 10912
rect 2996 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3162 10912
rect 2846 10847 3162 10848
rect 5846 10912 6162 10913
rect 5846 10848 5852 10912
rect 5916 10848 5932 10912
rect 5996 10848 6012 10912
rect 6076 10848 6092 10912
rect 6156 10848 6162 10912
rect 5846 10847 6162 10848
rect 8846 10912 9162 10913
rect 8846 10848 8852 10912
rect 8916 10848 8932 10912
rect 8996 10848 9012 10912
rect 9076 10848 9092 10912
rect 9156 10848 9162 10912
rect 8846 10847 9162 10848
rect 11846 10912 12162 10913
rect 11846 10848 11852 10912
rect 11916 10848 11932 10912
rect 11996 10848 12012 10912
rect 12076 10848 12092 10912
rect 12156 10848 12162 10912
rect 11846 10847 12162 10848
rect 14846 10912 15162 10913
rect 14846 10848 14852 10912
rect 14916 10848 14932 10912
rect 14996 10848 15012 10912
rect 15076 10848 15092 10912
rect 15156 10848 15162 10912
rect 14846 10847 15162 10848
rect 17846 10912 18162 10913
rect 17846 10848 17852 10912
rect 17916 10848 17932 10912
rect 17996 10848 18012 10912
rect 18076 10848 18092 10912
rect 18156 10848 18162 10912
rect 17846 10847 18162 10848
rect 20846 10912 21162 10913
rect 20846 10848 20852 10912
rect 20916 10848 20932 10912
rect 20996 10848 21012 10912
rect 21076 10848 21092 10912
rect 21156 10848 21162 10912
rect 20846 10847 21162 10848
rect 23846 10912 24162 10913
rect 23846 10848 23852 10912
rect 23916 10848 23932 10912
rect 23996 10848 24012 10912
rect 24076 10848 24092 10912
rect 24156 10848 24162 10912
rect 23846 10847 24162 10848
rect 6177 10706 6243 10709
rect 8201 10706 8267 10709
rect 6177 10704 8267 10706
rect 6177 10648 6182 10704
rect 6238 10648 8206 10704
rect 8262 10648 8267 10704
rect 6177 10646 8267 10648
rect 6177 10643 6243 10646
rect 8201 10643 8267 10646
rect 23289 10706 23355 10709
rect 24350 10706 24410 10918
rect 24780 10888 25180 10918
rect 23289 10704 24410 10706
rect 23289 10648 23294 10704
rect 23350 10648 24410 10704
rect 23289 10646 24410 10648
rect 23289 10643 23355 10646
rect 1853 10570 1919 10573
rect 982 10568 1919 10570
rect 982 10512 1858 10568
rect 1914 10512 1919 10568
rect 982 10510 1919 10512
rect 0 10298 400 10328
rect 982 10298 1042 10510
rect 1853 10507 1919 10510
rect 1346 10368 1662 10369
rect 1346 10304 1352 10368
rect 1416 10304 1432 10368
rect 1496 10304 1512 10368
rect 1576 10304 1592 10368
rect 1656 10304 1662 10368
rect 1346 10303 1662 10304
rect 4346 10368 4662 10369
rect 4346 10304 4352 10368
rect 4416 10304 4432 10368
rect 4496 10304 4512 10368
rect 4576 10304 4592 10368
rect 4656 10304 4662 10368
rect 4346 10303 4662 10304
rect 7346 10368 7662 10369
rect 7346 10304 7352 10368
rect 7416 10304 7432 10368
rect 7496 10304 7512 10368
rect 7576 10304 7592 10368
rect 7656 10304 7662 10368
rect 7346 10303 7662 10304
rect 10346 10368 10662 10369
rect 10346 10304 10352 10368
rect 10416 10304 10432 10368
rect 10496 10304 10512 10368
rect 10576 10304 10592 10368
rect 10656 10304 10662 10368
rect 10346 10303 10662 10304
rect 13346 10368 13662 10369
rect 13346 10304 13352 10368
rect 13416 10304 13432 10368
rect 13496 10304 13512 10368
rect 13576 10304 13592 10368
rect 13656 10304 13662 10368
rect 13346 10303 13662 10304
rect 16346 10368 16662 10369
rect 16346 10304 16352 10368
rect 16416 10304 16432 10368
rect 16496 10304 16512 10368
rect 16576 10304 16592 10368
rect 16656 10304 16662 10368
rect 16346 10303 16662 10304
rect 19346 10368 19662 10369
rect 19346 10304 19352 10368
rect 19416 10304 19432 10368
rect 19496 10304 19512 10368
rect 19576 10304 19592 10368
rect 19656 10304 19662 10368
rect 19346 10303 19662 10304
rect 22346 10368 22662 10369
rect 22346 10304 22352 10368
rect 22416 10304 22432 10368
rect 22496 10304 22512 10368
rect 22576 10304 22592 10368
rect 22656 10304 22662 10368
rect 22346 10303 22662 10304
rect 0 10238 1042 10298
rect 23381 10298 23447 10301
rect 24780 10298 25180 10328
rect 23381 10296 25180 10298
rect 23381 10240 23386 10296
rect 23442 10240 25180 10296
rect 23381 10238 25180 10240
rect 0 10208 400 10238
rect 23381 10235 23447 10238
rect 24780 10208 25180 10238
rect 2846 9824 3162 9825
rect 2846 9760 2852 9824
rect 2916 9760 2932 9824
rect 2996 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3162 9824
rect 2846 9759 3162 9760
rect 5846 9824 6162 9825
rect 5846 9760 5852 9824
rect 5916 9760 5932 9824
rect 5996 9760 6012 9824
rect 6076 9760 6092 9824
rect 6156 9760 6162 9824
rect 5846 9759 6162 9760
rect 8846 9824 9162 9825
rect 8846 9760 8852 9824
rect 8916 9760 8932 9824
rect 8996 9760 9012 9824
rect 9076 9760 9092 9824
rect 9156 9760 9162 9824
rect 8846 9759 9162 9760
rect 11846 9824 12162 9825
rect 11846 9760 11852 9824
rect 11916 9760 11932 9824
rect 11996 9760 12012 9824
rect 12076 9760 12092 9824
rect 12156 9760 12162 9824
rect 11846 9759 12162 9760
rect 14846 9824 15162 9825
rect 14846 9760 14852 9824
rect 14916 9760 14932 9824
rect 14996 9760 15012 9824
rect 15076 9760 15092 9824
rect 15156 9760 15162 9824
rect 14846 9759 15162 9760
rect 17846 9824 18162 9825
rect 17846 9760 17852 9824
rect 17916 9760 17932 9824
rect 17996 9760 18012 9824
rect 18076 9760 18092 9824
rect 18156 9760 18162 9824
rect 17846 9759 18162 9760
rect 20846 9824 21162 9825
rect 20846 9760 20852 9824
rect 20916 9760 20932 9824
rect 20996 9760 21012 9824
rect 21076 9760 21092 9824
rect 21156 9760 21162 9824
rect 20846 9759 21162 9760
rect 23846 9824 24162 9825
rect 23846 9760 23852 9824
rect 23916 9760 23932 9824
rect 23996 9760 24012 9824
rect 24076 9760 24092 9824
rect 24156 9760 24162 9824
rect 23846 9759 24162 9760
rect 0 9621 400 9648
rect 0 9616 447 9621
rect 0 9560 386 9616
rect 442 9560 447 9616
rect 0 9555 447 9560
rect 22829 9618 22895 9621
rect 24780 9618 25180 9648
rect 22829 9616 25180 9618
rect 22829 9560 22834 9616
rect 22890 9560 25180 9616
rect 22829 9558 25180 9560
rect 22829 9555 22895 9558
rect 0 9528 400 9555
rect 24780 9528 25180 9558
rect 1346 9280 1662 9281
rect 1346 9216 1352 9280
rect 1416 9216 1432 9280
rect 1496 9216 1512 9280
rect 1576 9216 1592 9280
rect 1656 9216 1662 9280
rect 1346 9215 1662 9216
rect 4346 9280 4662 9281
rect 4346 9216 4352 9280
rect 4416 9216 4432 9280
rect 4496 9216 4512 9280
rect 4576 9216 4592 9280
rect 4656 9216 4662 9280
rect 4346 9215 4662 9216
rect 7346 9280 7662 9281
rect 7346 9216 7352 9280
rect 7416 9216 7432 9280
rect 7496 9216 7512 9280
rect 7576 9216 7592 9280
rect 7656 9216 7662 9280
rect 7346 9215 7662 9216
rect 10346 9280 10662 9281
rect 10346 9216 10352 9280
rect 10416 9216 10432 9280
rect 10496 9216 10512 9280
rect 10576 9216 10592 9280
rect 10656 9216 10662 9280
rect 10346 9215 10662 9216
rect 13346 9280 13662 9281
rect 13346 9216 13352 9280
rect 13416 9216 13432 9280
rect 13496 9216 13512 9280
rect 13576 9216 13592 9280
rect 13656 9216 13662 9280
rect 13346 9215 13662 9216
rect 16346 9280 16662 9281
rect 16346 9216 16352 9280
rect 16416 9216 16432 9280
rect 16496 9216 16512 9280
rect 16576 9216 16592 9280
rect 16656 9216 16662 9280
rect 16346 9215 16662 9216
rect 19346 9280 19662 9281
rect 19346 9216 19352 9280
rect 19416 9216 19432 9280
rect 19496 9216 19512 9280
rect 19576 9216 19592 9280
rect 19656 9216 19662 9280
rect 19346 9215 19662 9216
rect 22346 9280 22662 9281
rect 22346 9216 22352 9280
rect 22416 9216 22432 9280
rect 22496 9216 22512 9280
rect 22576 9216 22592 9280
rect 22656 9216 22662 9280
rect 22346 9215 22662 9216
rect 0 8941 400 8968
rect 0 8936 447 8941
rect 0 8880 386 8936
rect 442 8880 447 8936
rect 0 8875 447 8880
rect 23381 8938 23447 8941
rect 24780 8938 25180 8968
rect 23381 8936 25180 8938
rect 23381 8880 23386 8936
rect 23442 8880 25180 8936
rect 23381 8878 25180 8880
rect 23381 8875 23447 8878
rect 0 8848 400 8875
rect 24780 8848 25180 8878
rect 2846 8736 3162 8737
rect 2846 8672 2852 8736
rect 2916 8672 2932 8736
rect 2996 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3162 8736
rect 2846 8671 3162 8672
rect 5846 8736 6162 8737
rect 5846 8672 5852 8736
rect 5916 8672 5932 8736
rect 5996 8672 6012 8736
rect 6076 8672 6092 8736
rect 6156 8672 6162 8736
rect 5846 8671 6162 8672
rect 8846 8736 9162 8737
rect 8846 8672 8852 8736
rect 8916 8672 8932 8736
rect 8996 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9162 8736
rect 8846 8671 9162 8672
rect 11846 8736 12162 8737
rect 11846 8672 11852 8736
rect 11916 8672 11932 8736
rect 11996 8672 12012 8736
rect 12076 8672 12092 8736
rect 12156 8672 12162 8736
rect 11846 8671 12162 8672
rect 14846 8736 15162 8737
rect 14846 8672 14852 8736
rect 14916 8672 14932 8736
rect 14996 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15162 8736
rect 14846 8671 15162 8672
rect 17846 8736 18162 8737
rect 17846 8672 17852 8736
rect 17916 8672 17932 8736
rect 17996 8672 18012 8736
rect 18076 8672 18092 8736
rect 18156 8672 18162 8736
rect 17846 8671 18162 8672
rect 20846 8736 21162 8737
rect 20846 8672 20852 8736
rect 20916 8672 20932 8736
rect 20996 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21162 8736
rect 20846 8671 21162 8672
rect 23846 8736 24162 8737
rect 23846 8672 23852 8736
rect 23916 8672 23932 8736
rect 23996 8672 24012 8736
rect 24076 8672 24092 8736
rect 24156 8672 24162 8736
rect 23846 8671 24162 8672
rect 14365 8394 14431 8397
rect 20621 8394 20687 8397
rect 14365 8392 20687 8394
rect 14365 8336 14370 8392
rect 14426 8336 20626 8392
rect 20682 8336 20687 8392
rect 14365 8334 20687 8336
rect 14365 8331 14431 8334
rect 0 8258 400 8288
rect 1209 8258 1275 8261
rect 0 8256 1275 8258
rect 0 8200 1214 8256
rect 1270 8200 1275 8256
rect 0 8198 1275 8200
rect 0 8168 400 8198
rect 1209 8195 1275 8198
rect 15193 8258 15259 8261
rect 15334 8258 15394 8334
rect 20621 8331 20687 8334
rect 15193 8256 15394 8258
rect 15193 8200 15198 8256
rect 15254 8200 15394 8256
rect 15193 8198 15394 8200
rect 15193 8195 15259 8198
rect 1346 8192 1662 8193
rect 1346 8128 1352 8192
rect 1416 8128 1432 8192
rect 1496 8128 1512 8192
rect 1576 8128 1592 8192
rect 1656 8128 1662 8192
rect 1346 8127 1662 8128
rect 4346 8192 4662 8193
rect 4346 8128 4352 8192
rect 4416 8128 4432 8192
rect 4496 8128 4512 8192
rect 4576 8128 4592 8192
rect 4656 8128 4662 8192
rect 4346 8127 4662 8128
rect 7346 8192 7662 8193
rect 7346 8128 7352 8192
rect 7416 8128 7432 8192
rect 7496 8128 7512 8192
rect 7576 8128 7592 8192
rect 7656 8128 7662 8192
rect 7346 8127 7662 8128
rect 10346 8192 10662 8193
rect 10346 8128 10352 8192
rect 10416 8128 10432 8192
rect 10496 8128 10512 8192
rect 10576 8128 10592 8192
rect 10656 8128 10662 8192
rect 10346 8127 10662 8128
rect 13346 8192 13662 8193
rect 13346 8128 13352 8192
rect 13416 8128 13432 8192
rect 13496 8128 13512 8192
rect 13576 8128 13592 8192
rect 13656 8128 13662 8192
rect 13346 8127 13662 8128
rect 16346 8192 16662 8193
rect 16346 8128 16352 8192
rect 16416 8128 16432 8192
rect 16496 8128 16512 8192
rect 16576 8128 16592 8192
rect 16656 8128 16662 8192
rect 16346 8127 16662 8128
rect 19346 8192 19662 8193
rect 19346 8128 19352 8192
rect 19416 8128 19432 8192
rect 19496 8128 19512 8192
rect 19576 8128 19592 8192
rect 19656 8128 19662 8192
rect 19346 8127 19662 8128
rect 22346 8192 22662 8193
rect 22346 8128 22352 8192
rect 22416 8128 22432 8192
rect 22496 8128 22512 8192
rect 22576 8128 22592 8192
rect 22656 8128 22662 8192
rect 22346 8127 22662 8128
rect 2846 7648 3162 7649
rect 2846 7584 2852 7648
rect 2916 7584 2932 7648
rect 2996 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3162 7648
rect 2846 7583 3162 7584
rect 5846 7648 6162 7649
rect 5846 7584 5852 7648
rect 5916 7584 5932 7648
rect 5996 7584 6012 7648
rect 6076 7584 6092 7648
rect 6156 7584 6162 7648
rect 5846 7583 6162 7584
rect 8846 7648 9162 7649
rect 8846 7584 8852 7648
rect 8916 7584 8932 7648
rect 8996 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9162 7648
rect 8846 7583 9162 7584
rect 11846 7648 12162 7649
rect 11846 7584 11852 7648
rect 11916 7584 11932 7648
rect 11996 7584 12012 7648
rect 12076 7584 12092 7648
rect 12156 7584 12162 7648
rect 11846 7583 12162 7584
rect 14846 7648 15162 7649
rect 14846 7584 14852 7648
rect 14916 7584 14932 7648
rect 14996 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15162 7648
rect 14846 7583 15162 7584
rect 17846 7648 18162 7649
rect 17846 7584 17852 7648
rect 17916 7584 17932 7648
rect 17996 7584 18012 7648
rect 18076 7584 18092 7648
rect 18156 7584 18162 7648
rect 17846 7583 18162 7584
rect 20846 7648 21162 7649
rect 20846 7584 20852 7648
rect 20916 7584 20932 7648
rect 20996 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21162 7648
rect 20846 7583 21162 7584
rect 23846 7648 24162 7649
rect 23846 7584 23852 7648
rect 23916 7584 23932 7648
rect 23996 7584 24012 7648
rect 24076 7584 24092 7648
rect 24156 7584 24162 7648
rect 23846 7583 24162 7584
rect 1346 7104 1662 7105
rect 1346 7040 1352 7104
rect 1416 7040 1432 7104
rect 1496 7040 1512 7104
rect 1576 7040 1592 7104
rect 1656 7040 1662 7104
rect 1346 7039 1662 7040
rect 4346 7104 4662 7105
rect 4346 7040 4352 7104
rect 4416 7040 4432 7104
rect 4496 7040 4512 7104
rect 4576 7040 4592 7104
rect 4656 7040 4662 7104
rect 4346 7039 4662 7040
rect 7346 7104 7662 7105
rect 7346 7040 7352 7104
rect 7416 7040 7432 7104
rect 7496 7040 7512 7104
rect 7576 7040 7592 7104
rect 7656 7040 7662 7104
rect 7346 7039 7662 7040
rect 10346 7104 10662 7105
rect 10346 7040 10352 7104
rect 10416 7040 10432 7104
rect 10496 7040 10512 7104
rect 10576 7040 10592 7104
rect 10656 7040 10662 7104
rect 10346 7039 10662 7040
rect 13346 7104 13662 7105
rect 13346 7040 13352 7104
rect 13416 7040 13432 7104
rect 13496 7040 13512 7104
rect 13576 7040 13592 7104
rect 13656 7040 13662 7104
rect 13346 7039 13662 7040
rect 16346 7104 16662 7105
rect 16346 7040 16352 7104
rect 16416 7040 16432 7104
rect 16496 7040 16512 7104
rect 16576 7040 16592 7104
rect 16656 7040 16662 7104
rect 16346 7039 16662 7040
rect 19346 7104 19662 7105
rect 19346 7040 19352 7104
rect 19416 7040 19432 7104
rect 19496 7040 19512 7104
rect 19576 7040 19592 7104
rect 19656 7040 19662 7104
rect 19346 7039 19662 7040
rect 22346 7104 22662 7105
rect 22346 7040 22352 7104
rect 22416 7040 22432 7104
rect 22496 7040 22512 7104
rect 22576 7040 22592 7104
rect 22656 7040 22662 7104
rect 22346 7039 22662 7040
rect 23381 6898 23447 6901
rect 24780 6898 25180 6928
rect 23381 6896 25180 6898
rect 23381 6840 23386 6896
rect 23442 6840 25180 6896
rect 23381 6838 25180 6840
rect 23381 6835 23447 6838
rect 24780 6808 25180 6838
rect 2846 6560 3162 6561
rect 2846 6496 2852 6560
rect 2916 6496 2932 6560
rect 2996 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3162 6560
rect 2846 6495 3162 6496
rect 5846 6560 6162 6561
rect 5846 6496 5852 6560
rect 5916 6496 5932 6560
rect 5996 6496 6012 6560
rect 6076 6496 6092 6560
rect 6156 6496 6162 6560
rect 5846 6495 6162 6496
rect 8846 6560 9162 6561
rect 8846 6496 8852 6560
rect 8916 6496 8932 6560
rect 8996 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9162 6560
rect 8846 6495 9162 6496
rect 11846 6560 12162 6561
rect 11846 6496 11852 6560
rect 11916 6496 11932 6560
rect 11996 6496 12012 6560
rect 12076 6496 12092 6560
rect 12156 6496 12162 6560
rect 11846 6495 12162 6496
rect 14846 6560 15162 6561
rect 14846 6496 14852 6560
rect 14916 6496 14932 6560
rect 14996 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15162 6560
rect 14846 6495 15162 6496
rect 17846 6560 18162 6561
rect 17846 6496 17852 6560
rect 17916 6496 17932 6560
rect 17996 6496 18012 6560
rect 18076 6496 18092 6560
rect 18156 6496 18162 6560
rect 17846 6495 18162 6496
rect 20846 6560 21162 6561
rect 20846 6496 20852 6560
rect 20916 6496 20932 6560
rect 20996 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21162 6560
rect 20846 6495 21162 6496
rect 23846 6560 24162 6561
rect 23846 6496 23852 6560
rect 23916 6496 23932 6560
rect 23996 6496 24012 6560
rect 24076 6496 24092 6560
rect 24156 6496 24162 6560
rect 23846 6495 24162 6496
rect 23657 6218 23723 6221
rect 24780 6218 25180 6248
rect 23657 6216 25180 6218
rect 23657 6160 23662 6216
rect 23718 6160 25180 6216
rect 23657 6158 25180 6160
rect 23657 6155 23723 6158
rect 24780 6128 25180 6158
rect 1346 6016 1662 6017
rect 1346 5952 1352 6016
rect 1416 5952 1432 6016
rect 1496 5952 1512 6016
rect 1576 5952 1592 6016
rect 1656 5952 1662 6016
rect 1346 5951 1662 5952
rect 4346 6016 4662 6017
rect 4346 5952 4352 6016
rect 4416 5952 4432 6016
rect 4496 5952 4512 6016
rect 4576 5952 4592 6016
rect 4656 5952 4662 6016
rect 4346 5951 4662 5952
rect 7346 6016 7662 6017
rect 7346 5952 7352 6016
rect 7416 5952 7432 6016
rect 7496 5952 7512 6016
rect 7576 5952 7592 6016
rect 7656 5952 7662 6016
rect 7346 5951 7662 5952
rect 10346 6016 10662 6017
rect 10346 5952 10352 6016
rect 10416 5952 10432 6016
rect 10496 5952 10512 6016
rect 10576 5952 10592 6016
rect 10656 5952 10662 6016
rect 10346 5951 10662 5952
rect 13346 6016 13662 6017
rect 13346 5952 13352 6016
rect 13416 5952 13432 6016
rect 13496 5952 13512 6016
rect 13576 5952 13592 6016
rect 13656 5952 13662 6016
rect 13346 5951 13662 5952
rect 16346 6016 16662 6017
rect 16346 5952 16352 6016
rect 16416 5952 16432 6016
rect 16496 5952 16512 6016
rect 16576 5952 16592 6016
rect 16656 5952 16662 6016
rect 16346 5951 16662 5952
rect 19346 6016 19662 6017
rect 19346 5952 19352 6016
rect 19416 5952 19432 6016
rect 19496 5952 19512 6016
rect 19576 5952 19592 6016
rect 19656 5952 19662 6016
rect 19346 5951 19662 5952
rect 22346 6016 22662 6017
rect 22346 5952 22352 6016
rect 22416 5952 22432 6016
rect 22496 5952 22512 6016
rect 22576 5952 22592 6016
rect 22656 5952 22662 6016
rect 22346 5951 22662 5952
rect 2846 5472 3162 5473
rect 2846 5408 2852 5472
rect 2916 5408 2932 5472
rect 2996 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3162 5472
rect 2846 5407 3162 5408
rect 5846 5472 6162 5473
rect 5846 5408 5852 5472
rect 5916 5408 5932 5472
rect 5996 5408 6012 5472
rect 6076 5408 6092 5472
rect 6156 5408 6162 5472
rect 5846 5407 6162 5408
rect 8846 5472 9162 5473
rect 8846 5408 8852 5472
rect 8916 5408 8932 5472
rect 8996 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9162 5472
rect 8846 5407 9162 5408
rect 11846 5472 12162 5473
rect 11846 5408 11852 5472
rect 11916 5408 11932 5472
rect 11996 5408 12012 5472
rect 12076 5408 12092 5472
rect 12156 5408 12162 5472
rect 11846 5407 12162 5408
rect 14846 5472 15162 5473
rect 14846 5408 14852 5472
rect 14916 5408 14932 5472
rect 14996 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15162 5472
rect 14846 5407 15162 5408
rect 17846 5472 18162 5473
rect 17846 5408 17852 5472
rect 17916 5408 17932 5472
rect 17996 5408 18012 5472
rect 18076 5408 18092 5472
rect 18156 5408 18162 5472
rect 17846 5407 18162 5408
rect 20846 5472 21162 5473
rect 20846 5408 20852 5472
rect 20916 5408 20932 5472
rect 20996 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21162 5472
rect 20846 5407 21162 5408
rect 23846 5472 24162 5473
rect 23846 5408 23852 5472
rect 23916 5408 23932 5472
rect 23996 5408 24012 5472
rect 24076 5408 24092 5472
rect 24156 5408 24162 5472
rect 23846 5407 24162 5408
rect 1346 4928 1662 4929
rect 1346 4864 1352 4928
rect 1416 4864 1432 4928
rect 1496 4864 1512 4928
rect 1576 4864 1592 4928
rect 1656 4864 1662 4928
rect 1346 4863 1662 4864
rect 4346 4928 4662 4929
rect 4346 4864 4352 4928
rect 4416 4864 4432 4928
rect 4496 4864 4512 4928
rect 4576 4864 4592 4928
rect 4656 4864 4662 4928
rect 4346 4863 4662 4864
rect 7346 4928 7662 4929
rect 7346 4864 7352 4928
rect 7416 4864 7432 4928
rect 7496 4864 7512 4928
rect 7576 4864 7592 4928
rect 7656 4864 7662 4928
rect 7346 4863 7662 4864
rect 10346 4928 10662 4929
rect 10346 4864 10352 4928
rect 10416 4864 10432 4928
rect 10496 4864 10512 4928
rect 10576 4864 10592 4928
rect 10656 4864 10662 4928
rect 10346 4863 10662 4864
rect 13346 4928 13662 4929
rect 13346 4864 13352 4928
rect 13416 4864 13432 4928
rect 13496 4864 13512 4928
rect 13576 4864 13592 4928
rect 13656 4864 13662 4928
rect 13346 4863 13662 4864
rect 16346 4928 16662 4929
rect 16346 4864 16352 4928
rect 16416 4864 16432 4928
rect 16496 4864 16512 4928
rect 16576 4864 16592 4928
rect 16656 4864 16662 4928
rect 16346 4863 16662 4864
rect 19346 4928 19662 4929
rect 19346 4864 19352 4928
rect 19416 4864 19432 4928
rect 19496 4864 19512 4928
rect 19576 4864 19592 4928
rect 19656 4864 19662 4928
rect 19346 4863 19662 4864
rect 22346 4928 22662 4929
rect 22346 4864 22352 4928
rect 22416 4864 22432 4928
rect 22496 4864 22512 4928
rect 22576 4864 22592 4928
rect 22656 4864 22662 4928
rect 22346 4863 22662 4864
rect 2846 4384 3162 4385
rect 2846 4320 2852 4384
rect 2916 4320 2932 4384
rect 2996 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3162 4384
rect 2846 4319 3162 4320
rect 5846 4384 6162 4385
rect 5846 4320 5852 4384
rect 5916 4320 5932 4384
rect 5996 4320 6012 4384
rect 6076 4320 6092 4384
rect 6156 4320 6162 4384
rect 5846 4319 6162 4320
rect 8846 4384 9162 4385
rect 8846 4320 8852 4384
rect 8916 4320 8932 4384
rect 8996 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9162 4384
rect 8846 4319 9162 4320
rect 11846 4384 12162 4385
rect 11846 4320 11852 4384
rect 11916 4320 11932 4384
rect 11996 4320 12012 4384
rect 12076 4320 12092 4384
rect 12156 4320 12162 4384
rect 11846 4319 12162 4320
rect 14846 4384 15162 4385
rect 14846 4320 14852 4384
rect 14916 4320 14932 4384
rect 14996 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15162 4384
rect 14846 4319 15162 4320
rect 17846 4384 18162 4385
rect 17846 4320 17852 4384
rect 17916 4320 17932 4384
rect 17996 4320 18012 4384
rect 18076 4320 18092 4384
rect 18156 4320 18162 4384
rect 17846 4319 18162 4320
rect 20846 4384 21162 4385
rect 20846 4320 20852 4384
rect 20916 4320 20932 4384
rect 20996 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21162 4384
rect 20846 4319 21162 4320
rect 23846 4384 24162 4385
rect 23846 4320 23852 4384
rect 23916 4320 23932 4384
rect 23996 4320 24012 4384
rect 24076 4320 24092 4384
rect 24156 4320 24162 4384
rect 23846 4319 24162 4320
rect 1346 3840 1662 3841
rect 1346 3776 1352 3840
rect 1416 3776 1432 3840
rect 1496 3776 1512 3840
rect 1576 3776 1592 3840
rect 1656 3776 1662 3840
rect 1346 3775 1662 3776
rect 4346 3840 4662 3841
rect 4346 3776 4352 3840
rect 4416 3776 4432 3840
rect 4496 3776 4512 3840
rect 4576 3776 4592 3840
rect 4656 3776 4662 3840
rect 4346 3775 4662 3776
rect 7346 3840 7662 3841
rect 7346 3776 7352 3840
rect 7416 3776 7432 3840
rect 7496 3776 7512 3840
rect 7576 3776 7592 3840
rect 7656 3776 7662 3840
rect 7346 3775 7662 3776
rect 10346 3840 10662 3841
rect 10346 3776 10352 3840
rect 10416 3776 10432 3840
rect 10496 3776 10512 3840
rect 10576 3776 10592 3840
rect 10656 3776 10662 3840
rect 10346 3775 10662 3776
rect 13346 3840 13662 3841
rect 13346 3776 13352 3840
rect 13416 3776 13432 3840
rect 13496 3776 13512 3840
rect 13576 3776 13592 3840
rect 13656 3776 13662 3840
rect 13346 3775 13662 3776
rect 16346 3840 16662 3841
rect 16346 3776 16352 3840
rect 16416 3776 16432 3840
rect 16496 3776 16512 3840
rect 16576 3776 16592 3840
rect 16656 3776 16662 3840
rect 16346 3775 16662 3776
rect 19346 3840 19662 3841
rect 19346 3776 19352 3840
rect 19416 3776 19432 3840
rect 19496 3776 19512 3840
rect 19576 3776 19592 3840
rect 19656 3776 19662 3840
rect 19346 3775 19662 3776
rect 22346 3840 22662 3841
rect 22346 3776 22352 3840
rect 22416 3776 22432 3840
rect 22496 3776 22512 3840
rect 22576 3776 22592 3840
rect 22656 3776 22662 3840
rect 22346 3775 22662 3776
rect 14733 3498 14799 3501
rect 16205 3498 16271 3501
rect 14733 3496 16271 3498
rect 14733 3440 14738 3496
rect 14794 3440 16210 3496
rect 16266 3440 16271 3496
rect 14733 3438 16271 3440
rect 14733 3435 14799 3438
rect 16205 3435 16271 3438
rect 2846 3296 3162 3297
rect 2846 3232 2852 3296
rect 2916 3232 2932 3296
rect 2996 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3162 3296
rect 2846 3231 3162 3232
rect 5846 3296 6162 3297
rect 5846 3232 5852 3296
rect 5916 3232 5932 3296
rect 5996 3232 6012 3296
rect 6076 3232 6092 3296
rect 6156 3232 6162 3296
rect 5846 3231 6162 3232
rect 8846 3296 9162 3297
rect 8846 3232 8852 3296
rect 8916 3232 8932 3296
rect 8996 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9162 3296
rect 8846 3231 9162 3232
rect 11846 3296 12162 3297
rect 11846 3232 11852 3296
rect 11916 3232 11932 3296
rect 11996 3232 12012 3296
rect 12076 3232 12092 3296
rect 12156 3232 12162 3296
rect 11846 3231 12162 3232
rect 14846 3296 15162 3297
rect 14846 3232 14852 3296
rect 14916 3232 14932 3296
rect 14996 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15162 3296
rect 14846 3231 15162 3232
rect 17846 3296 18162 3297
rect 17846 3232 17852 3296
rect 17916 3232 17932 3296
rect 17996 3232 18012 3296
rect 18076 3232 18092 3296
rect 18156 3232 18162 3296
rect 17846 3231 18162 3232
rect 20846 3296 21162 3297
rect 20846 3232 20852 3296
rect 20916 3232 20932 3296
rect 20996 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21162 3296
rect 20846 3231 21162 3232
rect 23846 3296 24162 3297
rect 23846 3232 23852 3296
rect 23916 3232 23932 3296
rect 23996 3232 24012 3296
rect 24076 3232 24092 3296
rect 24156 3232 24162 3296
rect 23846 3231 24162 3232
rect 1346 2752 1662 2753
rect 1346 2688 1352 2752
rect 1416 2688 1432 2752
rect 1496 2688 1512 2752
rect 1576 2688 1592 2752
rect 1656 2688 1662 2752
rect 1346 2687 1662 2688
rect 4346 2752 4662 2753
rect 4346 2688 4352 2752
rect 4416 2688 4432 2752
rect 4496 2688 4512 2752
rect 4576 2688 4592 2752
rect 4656 2688 4662 2752
rect 4346 2687 4662 2688
rect 7346 2752 7662 2753
rect 7346 2688 7352 2752
rect 7416 2688 7432 2752
rect 7496 2688 7512 2752
rect 7576 2688 7592 2752
rect 7656 2688 7662 2752
rect 7346 2687 7662 2688
rect 10346 2752 10662 2753
rect 10346 2688 10352 2752
rect 10416 2688 10432 2752
rect 10496 2688 10512 2752
rect 10576 2688 10592 2752
rect 10656 2688 10662 2752
rect 10346 2687 10662 2688
rect 13346 2752 13662 2753
rect 13346 2688 13352 2752
rect 13416 2688 13432 2752
rect 13496 2688 13512 2752
rect 13576 2688 13592 2752
rect 13656 2688 13662 2752
rect 13346 2687 13662 2688
rect 16346 2752 16662 2753
rect 16346 2688 16352 2752
rect 16416 2688 16432 2752
rect 16496 2688 16512 2752
rect 16576 2688 16592 2752
rect 16656 2688 16662 2752
rect 16346 2687 16662 2688
rect 19346 2752 19662 2753
rect 19346 2688 19352 2752
rect 19416 2688 19432 2752
rect 19496 2688 19512 2752
rect 19576 2688 19592 2752
rect 19656 2688 19662 2752
rect 19346 2687 19662 2688
rect 22346 2752 22662 2753
rect 22346 2688 22352 2752
rect 22416 2688 22432 2752
rect 22496 2688 22512 2752
rect 22576 2688 22592 2752
rect 22656 2688 22662 2752
rect 22346 2687 22662 2688
rect 2846 2208 3162 2209
rect 2846 2144 2852 2208
rect 2916 2144 2932 2208
rect 2996 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3162 2208
rect 2846 2143 3162 2144
rect 5846 2208 6162 2209
rect 5846 2144 5852 2208
rect 5916 2144 5932 2208
rect 5996 2144 6012 2208
rect 6076 2144 6092 2208
rect 6156 2144 6162 2208
rect 5846 2143 6162 2144
rect 8846 2208 9162 2209
rect 8846 2144 8852 2208
rect 8916 2144 8932 2208
rect 8996 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9162 2208
rect 8846 2143 9162 2144
rect 11846 2208 12162 2209
rect 11846 2144 11852 2208
rect 11916 2144 11932 2208
rect 11996 2144 12012 2208
rect 12076 2144 12092 2208
rect 12156 2144 12162 2208
rect 11846 2143 12162 2144
rect 14846 2208 15162 2209
rect 14846 2144 14852 2208
rect 14916 2144 14932 2208
rect 14996 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15162 2208
rect 14846 2143 15162 2144
rect 17846 2208 18162 2209
rect 17846 2144 17852 2208
rect 17916 2144 17932 2208
rect 17996 2144 18012 2208
rect 18076 2144 18092 2208
rect 18156 2144 18162 2208
rect 17846 2143 18162 2144
rect 20846 2208 21162 2209
rect 20846 2144 20852 2208
rect 20916 2144 20932 2208
rect 20996 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21162 2208
rect 20846 2143 21162 2144
rect 23846 2208 24162 2209
rect 23846 2144 23852 2208
rect 23916 2144 23932 2208
rect 23996 2144 24012 2208
rect 24076 2144 24092 2208
rect 24156 2144 24162 2208
rect 23846 2143 24162 2144
<< via3 >>
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 2932 25052 2996 25056
rect 2932 24996 2936 25052
rect 2936 24996 2992 25052
rect 2992 24996 2996 25052
rect 2932 24992 2996 24996
rect 3012 25052 3076 25056
rect 3012 24996 3016 25052
rect 3016 24996 3072 25052
rect 3072 24996 3076 25052
rect 3012 24992 3076 24996
rect 3092 25052 3156 25056
rect 3092 24996 3096 25052
rect 3096 24996 3152 25052
rect 3152 24996 3156 25052
rect 3092 24992 3156 24996
rect 5852 25052 5916 25056
rect 5852 24996 5856 25052
rect 5856 24996 5912 25052
rect 5912 24996 5916 25052
rect 5852 24992 5916 24996
rect 5932 25052 5996 25056
rect 5932 24996 5936 25052
rect 5936 24996 5992 25052
rect 5992 24996 5996 25052
rect 5932 24992 5996 24996
rect 6012 25052 6076 25056
rect 6012 24996 6016 25052
rect 6016 24996 6072 25052
rect 6072 24996 6076 25052
rect 6012 24992 6076 24996
rect 6092 25052 6156 25056
rect 6092 24996 6096 25052
rect 6096 24996 6152 25052
rect 6152 24996 6156 25052
rect 6092 24992 6156 24996
rect 8852 25052 8916 25056
rect 8852 24996 8856 25052
rect 8856 24996 8912 25052
rect 8912 24996 8916 25052
rect 8852 24992 8916 24996
rect 8932 25052 8996 25056
rect 8932 24996 8936 25052
rect 8936 24996 8992 25052
rect 8992 24996 8996 25052
rect 8932 24992 8996 24996
rect 9012 25052 9076 25056
rect 9012 24996 9016 25052
rect 9016 24996 9072 25052
rect 9072 24996 9076 25052
rect 9012 24992 9076 24996
rect 9092 25052 9156 25056
rect 9092 24996 9096 25052
rect 9096 24996 9152 25052
rect 9152 24996 9156 25052
rect 9092 24992 9156 24996
rect 11852 25052 11916 25056
rect 11852 24996 11856 25052
rect 11856 24996 11912 25052
rect 11912 24996 11916 25052
rect 11852 24992 11916 24996
rect 11932 25052 11996 25056
rect 11932 24996 11936 25052
rect 11936 24996 11992 25052
rect 11992 24996 11996 25052
rect 11932 24992 11996 24996
rect 12012 25052 12076 25056
rect 12012 24996 12016 25052
rect 12016 24996 12072 25052
rect 12072 24996 12076 25052
rect 12012 24992 12076 24996
rect 12092 25052 12156 25056
rect 12092 24996 12096 25052
rect 12096 24996 12152 25052
rect 12152 24996 12156 25052
rect 12092 24992 12156 24996
rect 14852 25052 14916 25056
rect 14852 24996 14856 25052
rect 14856 24996 14912 25052
rect 14912 24996 14916 25052
rect 14852 24992 14916 24996
rect 14932 25052 14996 25056
rect 14932 24996 14936 25052
rect 14936 24996 14992 25052
rect 14992 24996 14996 25052
rect 14932 24992 14996 24996
rect 15012 25052 15076 25056
rect 15012 24996 15016 25052
rect 15016 24996 15072 25052
rect 15072 24996 15076 25052
rect 15012 24992 15076 24996
rect 15092 25052 15156 25056
rect 15092 24996 15096 25052
rect 15096 24996 15152 25052
rect 15152 24996 15156 25052
rect 15092 24992 15156 24996
rect 17852 25052 17916 25056
rect 17852 24996 17856 25052
rect 17856 24996 17912 25052
rect 17912 24996 17916 25052
rect 17852 24992 17916 24996
rect 17932 25052 17996 25056
rect 17932 24996 17936 25052
rect 17936 24996 17992 25052
rect 17992 24996 17996 25052
rect 17932 24992 17996 24996
rect 18012 25052 18076 25056
rect 18012 24996 18016 25052
rect 18016 24996 18072 25052
rect 18072 24996 18076 25052
rect 18012 24992 18076 24996
rect 18092 25052 18156 25056
rect 18092 24996 18096 25052
rect 18096 24996 18152 25052
rect 18152 24996 18156 25052
rect 18092 24992 18156 24996
rect 20852 25052 20916 25056
rect 20852 24996 20856 25052
rect 20856 24996 20912 25052
rect 20912 24996 20916 25052
rect 20852 24992 20916 24996
rect 20932 25052 20996 25056
rect 20932 24996 20936 25052
rect 20936 24996 20992 25052
rect 20992 24996 20996 25052
rect 20932 24992 20996 24996
rect 21012 25052 21076 25056
rect 21012 24996 21016 25052
rect 21016 24996 21072 25052
rect 21072 24996 21076 25052
rect 21012 24992 21076 24996
rect 21092 25052 21156 25056
rect 21092 24996 21096 25052
rect 21096 24996 21152 25052
rect 21152 24996 21156 25052
rect 21092 24992 21156 24996
rect 23852 25052 23916 25056
rect 23852 24996 23856 25052
rect 23856 24996 23912 25052
rect 23912 24996 23916 25052
rect 23852 24992 23916 24996
rect 23932 25052 23996 25056
rect 23932 24996 23936 25052
rect 23936 24996 23992 25052
rect 23992 24996 23996 25052
rect 23932 24992 23996 24996
rect 24012 25052 24076 25056
rect 24012 24996 24016 25052
rect 24016 24996 24072 25052
rect 24072 24996 24076 25052
rect 24012 24992 24076 24996
rect 24092 25052 24156 25056
rect 24092 24996 24096 25052
rect 24096 24996 24152 25052
rect 24152 24996 24156 25052
rect 24092 24992 24156 24996
rect 1352 24508 1416 24512
rect 1352 24452 1356 24508
rect 1356 24452 1412 24508
rect 1412 24452 1416 24508
rect 1352 24448 1416 24452
rect 1432 24508 1496 24512
rect 1432 24452 1436 24508
rect 1436 24452 1492 24508
rect 1492 24452 1496 24508
rect 1432 24448 1496 24452
rect 1512 24508 1576 24512
rect 1512 24452 1516 24508
rect 1516 24452 1572 24508
rect 1572 24452 1576 24508
rect 1512 24448 1576 24452
rect 1592 24508 1656 24512
rect 1592 24452 1596 24508
rect 1596 24452 1652 24508
rect 1652 24452 1656 24508
rect 1592 24448 1656 24452
rect 4352 24508 4416 24512
rect 4352 24452 4356 24508
rect 4356 24452 4412 24508
rect 4412 24452 4416 24508
rect 4352 24448 4416 24452
rect 4432 24508 4496 24512
rect 4432 24452 4436 24508
rect 4436 24452 4492 24508
rect 4492 24452 4496 24508
rect 4432 24448 4496 24452
rect 4512 24508 4576 24512
rect 4512 24452 4516 24508
rect 4516 24452 4572 24508
rect 4572 24452 4576 24508
rect 4512 24448 4576 24452
rect 4592 24508 4656 24512
rect 4592 24452 4596 24508
rect 4596 24452 4652 24508
rect 4652 24452 4656 24508
rect 4592 24448 4656 24452
rect 7352 24508 7416 24512
rect 7352 24452 7356 24508
rect 7356 24452 7412 24508
rect 7412 24452 7416 24508
rect 7352 24448 7416 24452
rect 7432 24508 7496 24512
rect 7432 24452 7436 24508
rect 7436 24452 7492 24508
rect 7492 24452 7496 24508
rect 7432 24448 7496 24452
rect 7512 24508 7576 24512
rect 7512 24452 7516 24508
rect 7516 24452 7572 24508
rect 7572 24452 7576 24508
rect 7512 24448 7576 24452
rect 7592 24508 7656 24512
rect 7592 24452 7596 24508
rect 7596 24452 7652 24508
rect 7652 24452 7656 24508
rect 7592 24448 7656 24452
rect 10352 24508 10416 24512
rect 10352 24452 10356 24508
rect 10356 24452 10412 24508
rect 10412 24452 10416 24508
rect 10352 24448 10416 24452
rect 10432 24508 10496 24512
rect 10432 24452 10436 24508
rect 10436 24452 10492 24508
rect 10492 24452 10496 24508
rect 10432 24448 10496 24452
rect 10512 24508 10576 24512
rect 10512 24452 10516 24508
rect 10516 24452 10572 24508
rect 10572 24452 10576 24508
rect 10512 24448 10576 24452
rect 10592 24508 10656 24512
rect 10592 24452 10596 24508
rect 10596 24452 10652 24508
rect 10652 24452 10656 24508
rect 10592 24448 10656 24452
rect 13352 24508 13416 24512
rect 13352 24452 13356 24508
rect 13356 24452 13412 24508
rect 13412 24452 13416 24508
rect 13352 24448 13416 24452
rect 13432 24508 13496 24512
rect 13432 24452 13436 24508
rect 13436 24452 13492 24508
rect 13492 24452 13496 24508
rect 13432 24448 13496 24452
rect 13512 24508 13576 24512
rect 13512 24452 13516 24508
rect 13516 24452 13572 24508
rect 13572 24452 13576 24508
rect 13512 24448 13576 24452
rect 13592 24508 13656 24512
rect 13592 24452 13596 24508
rect 13596 24452 13652 24508
rect 13652 24452 13656 24508
rect 13592 24448 13656 24452
rect 16352 24508 16416 24512
rect 16352 24452 16356 24508
rect 16356 24452 16412 24508
rect 16412 24452 16416 24508
rect 16352 24448 16416 24452
rect 16432 24508 16496 24512
rect 16432 24452 16436 24508
rect 16436 24452 16492 24508
rect 16492 24452 16496 24508
rect 16432 24448 16496 24452
rect 16512 24508 16576 24512
rect 16512 24452 16516 24508
rect 16516 24452 16572 24508
rect 16572 24452 16576 24508
rect 16512 24448 16576 24452
rect 16592 24508 16656 24512
rect 16592 24452 16596 24508
rect 16596 24452 16652 24508
rect 16652 24452 16656 24508
rect 16592 24448 16656 24452
rect 19352 24508 19416 24512
rect 19352 24452 19356 24508
rect 19356 24452 19412 24508
rect 19412 24452 19416 24508
rect 19352 24448 19416 24452
rect 19432 24508 19496 24512
rect 19432 24452 19436 24508
rect 19436 24452 19492 24508
rect 19492 24452 19496 24508
rect 19432 24448 19496 24452
rect 19512 24508 19576 24512
rect 19512 24452 19516 24508
rect 19516 24452 19572 24508
rect 19572 24452 19576 24508
rect 19512 24448 19576 24452
rect 19592 24508 19656 24512
rect 19592 24452 19596 24508
rect 19596 24452 19652 24508
rect 19652 24452 19656 24508
rect 19592 24448 19656 24452
rect 22352 24508 22416 24512
rect 22352 24452 22356 24508
rect 22356 24452 22412 24508
rect 22412 24452 22416 24508
rect 22352 24448 22416 24452
rect 22432 24508 22496 24512
rect 22432 24452 22436 24508
rect 22436 24452 22492 24508
rect 22492 24452 22496 24508
rect 22432 24448 22496 24452
rect 22512 24508 22576 24512
rect 22512 24452 22516 24508
rect 22516 24452 22572 24508
rect 22572 24452 22576 24508
rect 22512 24448 22576 24452
rect 22592 24508 22656 24512
rect 22592 24452 22596 24508
rect 22596 24452 22652 24508
rect 22652 24452 22656 24508
rect 22592 24448 22656 24452
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 2932 23964 2996 23968
rect 2932 23908 2936 23964
rect 2936 23908 2992 23964
rect 2992 23908 2996 23964
rect 2932 23904 2996 23908
rect 3012 23964 3076 23968
rect 3012 23908 3016 23964
rect 3016 23908 3072 23964
rect 3072 23908 3076 23964
rect 3012 23904 3076 23908
rect 3092 23964 3156 23968
rect 3092 23908 3096 23964
rect 3096 23908 3152 23964
rect 3152 23908 3156 23964
rect 3092 23904 3156 23908
rect 5852 23964 5916 23968
rect 5852 23908 5856 23964
rect 5856 23908 5912 23964
rect 5912 23908 5916 23964
rect 5852 23904 5916 23908
rect 5932 23964 5996 23968
rect 5932 23908 5936 23964
rect 5936 23908 5992 23964
rect 5992 23908 5996 23964
rect 5932 23904 5996 23908
rect 6012 23964 6076 23968
rect 6012 23908 6016 23964
rect 6016 23908 6072 23964
rect 6072 23908 6076 23964
rect 6012 23904 6076 23908
rect 6092 23964 6156 23968
rect 6092 23908 6096 23964
rect 6096 23908 6152 23964
rect 6152 23908 6156 23964
rect 6092 23904 6156 23908
rect 8852 23964 8916 23968
rect 8852 23908 8856 23964
rect 8856 23908 8912 23964
rect 8912 23908 8916 23964
rect 8852 23904 8916 23908
rect 8932 23964 8996 23968
rect 8932 23908 8936 23964
rect 8936 23908 8992 23964
rect 8992 23908 8996 23964
rect 8932 23904 8996 23908
rect 9012 23964 9076 23968
rect 9012 23908 9016 23964
rect 9016 23908 9072 23964
rect 9072 23908 9076 23964
rect 9012 23904 9076 23908
rect 9092 23964 9156 23968
rect 9092 23908 9096 23964
rect 9096 23908 9152 23964
rect 9152 23908 9156 23964
rect 9092 23904 9156 23908
rect 11852 23964 11916 23968
rect 11852 23908 11856 23964
rect 11856 23908 11912 23964
rect 11912 23908 11916 23964
rect 11852 23904 11916 23908
rect 11932 23964 11996 23968
rect 11932 23908 11936 23964
rect 11936 23908 11992 23964
rect 11992 23908 11996 23964
rect 11932 23904 11996 23908
rect 12012 23964 12076 23968
rect 12012 23908 12016 23964
rect 12016 23908 12072 23964
rect 12072 23908 12076 23964
rect 12012 23904 12076 23908
rect 12092 23964 12156 23968
rect 12092 23908 12096 23964
rect 12096 23908 12152 23964
rect 12152 23908 12156 23964
rect 12092 23904 12156 23908
rect 14852 23964 14916 23968
rect 14852 23908 14856 23964
rect 14856 23908 14912 23964
rect 14912 23908 14916 23964
rect 14852 23904 14916 23908
rect 14932 23964 14996 23968
rect 14932 23908 14936 23964
rect 14936 23908 14992 23964
rect 14992 23908 14996 23964
rect 14932 23904 14996 23908
rect 15012 23964 15076 23968
rect 15012 23908 15016 23964
rect 15016 23908 15072 23964
rect 15072 23908 15076 23964
rect 15012 23904 15076 23908
rect 15092 23964 15156 23968
rect 15092 23908 15096 23964
rect 15096 23908 15152 23964
rect 15152 23908 15156 23964
rect 15092 23904 15156 23908
rect 17852 23964 17916 23968
rect 17852 23908 17856 23964
rect 17856 23908 17912 23964
rect 17912 23908 17916 23964
rect 17852 23904 17916 23908
rect 17932 23964 17996 23968
rect 17932 23908 17936 23964
rect 17936 23908 17992 23964
rect 17992 23908 17996 23964
rect 17932 23904 17996 23908
rect 18012 23964 18076 23968
rect 18012 23908 18016 23964
rect 18016 23908 18072 23964
rect 18072 23908 18076 23964
rect 18012 23904 18076 23908
rect 18092 23964 18156 23968
rect 18092 23908 18096 23964
rect 18096 23908 18152 23964
rect 18152 23908 18156 23964
rect 18092 23904 18156 23908
rect 20852 23964 20916 23968
rect 20852 23908 20856 23964
rect 20856 23908 20912 23964
rect 20912 23908 20916 23964
rect 20852 23904 20916 23908
rect 20932 23964 20996 23968
rect 20932 23908 20936 23964
rect 20936 23908 20992 23964
rect 20992 23908 20996 23964
rect 20932 23904 20996 23908
rect 21012 23964 21076 23968
rect 21012 23908 21016 23964
rect 21016 23908 21072 23964
rect 21072 23908 21076 23964
rect 21012 23904 21076 23908
rect 21092 23964 21156 23968
rect 21092 23908 21096 23964
rect 21096 23908 21152 23964
rect 21152 23908 21156 23964
rect 21092 23904 21156 23908
rect 23852 23964 23916 23968
rect 23852 23908 23856 23964
rect 23856 23908 23912 23964
rect 23912 23908 23916 23964
rect 23852 23904 23916 23908
rect 23932 23964 23996 23968
rect 23932 23908 23936 23964
rect 23936 23908 23992 23964
rect 23992 23908 23996 23964
rect 23932 23904 23996 23908
rect 24012 23964 24076 23968
rect 24012 23908 24016 23964
rect 24016 23908 24072 23964
rect 24072 23908 24076 23964
rect 24012 23904 24076 23908
rect 24092 23964 24156 23968
rect 24092 23908 24096 23964
rect 24096 23908 24152 23964
rect 24152 23908 24156 23964
rect 24092 23904 24156 23908
rect 1352 23420 1416 23424
rect 1352 23364 1356 23420
rect 1356 23364 1412 23420
rect 1412 23364 1416 23420
rect 1352 23360 1416 23364
rect 1432 23420 1496 23424
rect 1432 23364 1436 23420
rect 1436 23364 1492 23420
rect 1492 23364 1496 23420
rect 1432 23360 1496 23364
rect 1512 23420 1576 23424
rect 1512 23364 1516 23420
rect 1516 23364 1572 23420
rect 1572 23364 1576 23420
rect 1512 23360 1576 23364
rect 1592 23420 1656 23424
rect 1592 23364 1596 23420
rect 1596 23364 1652 23420
rect 1652 23364 1656 23420
rect 1592 23360 1656 23364
rect 4352 23420 4416 23424
rect 4352 23364 4356 23420
rect 4356 23364 4412 23420
rect 4412 23364 4416 23420
rect 4352 23360 4416 23364
rect 4432 23420 4496 23424
rect 4432 23364 4436 23420
rect 4436 23364 4492 23420
rect 4492 23364 4496 23420
rect 4432 23360 4496 23364
rect 4512 23420 4576 23424
rect 4512 23364 4516 23420
rect 4516 23364 4572 23420
rect 4572 23364 4576 23420
rect 4512 23360 4576 23364
rect 4592 23420 4656 23424
rect 4592 23364 4596 23420
rect 4596 23364 4652 23420
rect 4652 23364 4656 23420
rect 4592 23360 4656 23364
rect 7352 23420 7416 23424
rect 7352 23364 7356 23420
rect 7356 23364 7412 23420
rect 7412 23364 7416 23420
rect 7352 23360 7416 23364
rect 7432 23420 7496 23424
rect 7432 23364 7436 23420
rect 7436 23364 7492 23420
rect 7492 23364 7496 23420
rect 7432 23360 7496 23364
rect 7512 23420 7576 23424
rect 7512 23364 7516 23420
rect 7516 23364 7572 23420
rect 7572 23364 7576 23420
rect 7512 23360 7576 23364
rect 7592 23420 7656 23424
rect 7592 23364 7596 23420
rect 7596 23364 7652 23420
rect 7652 23364 7656 23420
rect 7592 23360 7656 23364
rect 10352 23420 10416 23424
rect 10352 23364 10356 23420
rect 10356 23364 10412 23420
rect 10412 23364 10416 23420
rect 10352 23360 10416 23364
rect 10432 23420 10496 23424
rect 10432 23364 10436 23420
rect 10436 23364 10492 23420
rect 10492 23364 10496 23420
rect 10432 23360 10496 23364
rect 10512 23420 10576 23424
rect 10512 23364 10516 23420
rect 10516 23364 10572 23420
rect 10572 23364 10576 23420
rect 10512 23360 10576 23364
rect 10592 23420 10656 23424
rect 10592 23364 10596 23420
rect 10596 23364 10652 23420
rect 10652 23364 10656 23420
rect 10592 23360 10656 23364
rect 13352 23420 13416 23424
rect 13352 23364 13356 23420
rect 13356 23364 13412 23420
rect 13412 23364 13416 23420
rect 13352 23360 13416 23364
rect 13432 23420 13496 23424
rect 13432 23364 13436 23420
rect 13436 23364 13492 23420
rect 13492 23364 13496 23420
rect 13432 23360 13496 23364
rect 13512 23420 13576 23424
rect 13512 23364 13516 23420
rect 13516 23364 13572 23420
rect 13572 23364 13576 23420
rect 13512 23360 13576 23364
rect 13592 23420 13656 23424
rect 13592 23364 13596 23420
rect 13596 23364 13652 23420
rect 13652 23364 13656 23420
rect 13592 23360 13656 23364
rect 16352 23420 16416 23424
rect 16352 23364 16356 23420
rect 16356 23364 16412 23420
rect 16412 23364 16416 23420
rect 16352 23360 16416 23364
rect 16432 23420 16496 23424
rect 16432 23364 16436 23420
rect 16436 23364 16492 23420
rect 16492 23364 16496 23420
rect 16432 23360 16496 23364
rect 16512 23420 16576 23424
rect 16512 23364 16516 23420
rect 16516 23364 16572 23420
rect 16572 23364 16576 23420
rect 16512 23360 16576 23364
rect 16592 23420 16656 23424
rect 16592 23364 16596 23420
rect 16596 23364 16652 23420
rect 16652 23364 16656 23420
rect 16592 23360 16656 23364
rect 19352 23420 19416 23424
rect 19352 23364 19356 23420
rect 19356 23364 19412 23420
rect 19412 23364 19416 23420
rect 19352 23360 19416 23364
rect 19432 23420 19496 23424
rect 19432 23364 19436 23420
rect 19436 23364 19492 23420
rect 19492 23364 19496 23420
rect 19432 23360 19496 23364
rect 19512 23420 19576 23424
rect 19512 23364 19516 23420
rect 19516 23364 19572 23420
rect 19572 23364 19576 23420
rect 19512 23360 19576 23364
rect 19592 23420 19656 23424
rect 19592 23364 19596 23420
rect 19596 23364 19652 23420
rect 19652 23364 19656 23420
rect 19592 23360 19656 23364
rect 22352 23420 22416 23424
rect 22352 23364 22356 23420
rect 22356 23364 22412 23420
rect 22412 23364 22416 23420
rect 22352 23360 22416 23364
rect 22432 23420 22496 23424
rect 22432 23364 22436 23420
rect 22436 23364 22492 23420
rect 22492 23364 22496 23420
rect 22432 23360 22496 23364
rect 22512 23420 22576 23424
rect 22512 23364 22516 23420
rect 22516 23364 22572 23420
rect 22572 23364 22576 23420
rect 22512 23360 22576 23364
rect 22592 23420 22656 23424
rect 22592 23364 22596 23420
rect 22596 23364 22652 23420
rect 22652 23364 22656 23420
rect 22592 23360 22656 23364
rect 3372 23156 3436 23220
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 2932 22876 2996 22880
rect 2932 22820 2936 22876
rect 2936 22820 2992 22876
rect 2992 22820 2996 22876
rect 2932 22816 2996 22820
rect 3012 22876 3076 22880
rect 3012 22820 3016 22876
rect 3016 22820 3072 22876
rect 3072 22820 3076 22876
rect 3012 22816 3076 22820
rect 3092 22876 3156 22880
rect 3092 22820 3096 22876
rect 3096 22820 3152 22876
rect 3152 22820 3156 22876
rect 3092 22816 3156 22820
rect 5852 22876 5916 22880
rect 5852 22820 5856 22876
rect 5856 22820 5912 22876
rect 5912 22820 5916 22876
rect 5852 22816 5916 22820
rect 5932 22876 5996 22880
rect 5932 22820 5936 22876
rect 5936 22820 5992 22876
rect 5992 22820 5996 22876
rect 5932 22816 5996 22820
rect 6012 22876 6076 22880
rect 6012 22820 6016 22876
rect 6016 22820 6072 22876
rect 6072 22820 6076 22876
rect 6012 22816 6076 22820
rect 6092 22876 6156 22880
rect 6092 22820 6096 22876
rect 6096 22820 6152 22876
rect 6152 22820 6156 22876
rect 6092 22816 6156 22820
rect 8852 22876 8916 22880
rect 8852 22820 8856 22876
rect 8856 22820 8912 22876
rect 8912 22820 8916 22876
rect 8852 22816 8916 22820
rect 8932 22876 8996 22880
rect 8932 22820 8936 22876
rect 8936 22820 8992 22876
rect 8992 22820 8996 22876
rect 8932 22816 8996 22820
rect 9012 22876 9076 22880
rect 9012 22820 9016 22876
rect 9016 22820 9072 22876
rect 9072 22820 9076 22876
rect 9012 22816 9076 22820
rect 9092 22876 9156 22880
rect 9092 22820 9096 22876
rect 9096 22820 9152 22876
rect 9152 22820 9156 22876
rect 9092 22816 9156 22820
rect 11852 22876 11916 22880
rect 11852 22820 11856 22876
rect 11856 22820 11912 22876
rect 11912 22820 11916 22876
rect 11852 22816 11916 22820
rect 11932 22876 11996 22880
rect 11932 22820 11936 22876
rect 11936 22820 11992 22876
rect 11992 22820 11996 22876
rect 11932 22816 11996 22820
rect 12012 22876 12076 22880
rect 12012 22820 12016 22876
rect 12016 22820 12072 22876
rect 12072 22820 12076 22876
rect 12012 22816 12076 22820
rect 12092 22876 12156 22880
rect 12092 22820 12096 22876
rect 12096 22820 12152 22876
rect 12152 22820 12156 22876
rect 12092 22816 12156 22820
rect 14852 22876 14916 22880
rect 14852 22820 14856 22876
rect 14856 22820 14912 22876
rect 14912 22820 14916 22876
rect 14852 22816 14916 22820
rect 14932 22876 14996 22880
rect 14932 22820 14936 22876
rect 14936 22820 14992 22876
rect 14992 22820 14996 22876
rect 14932 22816 14996 22820
rect 15012 22876 15076 22880
rect 15012 22820 15016 22876
rect 15016 22820 15072 22876
rect 15072 22820 15076 22876
rect 15012 22816 15076 22820
rect 15092 22876 15156 22880
rect 15092 22820 15096 22876
rect 15096 22820 15152 22876
rect 15152 22820 15156 22876
rect 15092 22816 15156 22820
rect 17852 22876 17916 22880
rect 17852 22820 17856 22876
rect 17856 22820 17912 22876
rect 17912 22820 17916 22876
rect 17852 22816 17916 22820
rect 17932 22876 17996 22880
rect 17932 22820 17936 22876
rect 17936 22820 17992 22876
rect 17992 22820 17996 22876
rect 17932 22816 17996 22820
rect 18012 22876 18076 22880
rect 18012 22820 18016 22876
rect 18016 22820 18072 22876
rect 18072 22820 18076 22876
rect 18012 22816 18076 22820
rect 18092 22876 18156 22880
rect 18092 22820 18096 22876
rect 18096 22820 18152 22876
rect 18152 22820 18156 22876
rect 18092 22816 18156 22820
rect 20852 22876 20916 22880
rect 20852 22820 20856 22876
rect 20856 22820 20912 22876
rect 20912 22820 20916 22876
rect 20852 22816 20916 22820
rect 20932 22876 20996 22880
rect 20932 22820 20936 22876
rect 20936 22820 20992 22876
rect 20992 22820 20996 22876
rect 20932 22816 20996 22820
rect 21012 22876 21076 22880
rect 21012 22820 21016 22876
rect 21016 22820 21072 22876
rect 21072 22820 21076 22876
rect 21012 22816 21076 22820
rect 21092 22876 21156 22880
rect 21092 22820 21096 22876
rect 21096 22820 21152 22876
rect 21152 22820 21156 22876
rect 21092 22816 21156 22820
rect 23852 22876 23916 22880
rect 23852 22820 23856 22876
rect 23856 22820 23912 22876
rect 23912 22820 23916 22876
rect 23852 22816 23916 22820
rect 23932 22876 23996 22880
rect 23932 22820 23936 22876
rect 23936 22820 23992 22876
rect 23992 22820 23996 22876
rect 23932 22816 23996 22820
rect 24012 22876 24076 22880
rect 24012 22820 24016 22876
rect 24016 22820 24072 22876
rect 24072 22820 24076 22876
rect 24012 22816 24076 22820
rect 24092 22876 24156 22880
rect 24092 22820 24096 22876
rect 24096 22820 24152 22876
rect 24152 22820 24156 22876
rect 24092 22816 24156 22820
rect 1352 22332 1416 22336
rect 1352 22276 1356 22332
rect 1356 22276 1412 22332
rect 1412 22276 1416 22332
rect 1352 22272 1416 22276
rect 1432 22332 1496 22336
rect 1432 22276 1436 22332
rect 1436 22276 1492 22332
rect 1492 22276 1496 22332
rect 1432 22272 1496 22276
rect 1512 22332 1576 22336
rect 1512 22276 1516 22332
rect 1516 22276 1572 22332
rect 1572 22276 1576 22332
rect 1512 22272 1576 22276
rect 1592 22332 1656 22336
rect 1592 22276 1596 22332
rect 1596 22276 1652 22332
rect 1652 22276 1656 22332
rect 1592 22272 1656 22276
rect 4352 22332 4416 22336
rect 4352 22276 4356 22332
rect 4356 22276 4412 22332
rect 4412 22276 4416 22332
rect 4352 22272 4416 22276
rect 4432 22332 4496 22336
rect 4432 22276 4436 22332
rect 4436 22276 4492 22332
rect 4492 22276 4496 22332
rect 4432 22272 4496 22276
rect 4512 22332 4576 22336
rect 4512 22276 4516 22332
rect 4516 22276 4572 22332
rect 4572 22276 4576 22332
rect 4512 22272 4576 22276
rect 4592 22332 4656 22336
rect 4592 22276 4596 22332
rect 4596 22276 4652 22332
rect 4652 22276 4656 22332
rect 4592 22272 4656 22276
rect 7352 22332 7416 22336
rect 7352 22276 7356 22332
rect 7356 22276 7412 22332
rect 7412 22276 7416 22332
rect 7352 22272 7416 22276
rect 7432 22332 7496 22336
rect 7432 22276 7436 22332
rect 7436 22276 7492 22332
rect 7492 22276 7496 22332
rect 7432 22272 7496 22276
rect 7512 22332 7576 22336
rect 7512 22276 7516 22332
rect 7516 22276 7572 22332
rect 7572 22276 7576 22332
rect 7512 22272 7576 22276
rect 7592 22332 7656 22336
rect 7592 22276 7596 22332
rect 7596 22276 7652 22332
rect 7652 22276 7656 22332
rect 7592 22272 7656 22276
rect 10352 22332 10416 22336
rect 10352 22276 10356 22332
rect 10356 22276 10412 22332
rect 10412 22276 10416 22332
rect 10352 22272 10416 22276
rect 10432 22332 10496 22336
rect 10432 22276 10436 22332
rect 10436 22276 10492 22332
rect 10492 22276 10496 22332
rect 10432 22272 10496 22276
rect 10512 22332 10576 22336
rect 10512 22276 10516 22332
rect 10516 22276 10572 22332
rect 10572 22276 10576 22332
rect 10512 22272 10576 22276
rect 10592 22332 10656 22336
rect 10592 22276 10596 22332
rect 10596 22276 10652 22332
rect 10652 22276 10656 22332
rect 10592 22272 10656 22276
rect 13352 22332 13416 22336
rect 13352 22276 13356 22332
rect 13356 22276 13412 22332
rect 13412 22276 13416 22332
rect 13352 22272 13416 22276
rect 13432 22332 13496 22336
rect 13432 22276 13436 22332
rect 13436 22276 13492 22332
rect 13492 22276 13496 22332
rect 13432 22272 13496 22276
rect 13512 22332 13576 22336
rect 13512 22276 13516 22332
rect 13516 22276 13572 22332
rect 13572 22276 13576 22332
rect 13512 22272 13576 22276
rect 13592 22332 13656 22336
rect 13592 22276 13596 22332
rect 13596 22276 13652 22332
rect 13652 22276 13656 22332
rect 13592 22272 13656 22276
rect 16352 22332 16416 22336
rect 16352 22276 16356 22332
rect 16356 22276 16412 22332
rect 16412 22276 16416 22332
rect 16352 22272 16416 22276
rect 16432 22332 16496 22336
rect 16432 22276 16436 22332
rect 16436 22276 16492 22332
rect 16492 22276 16496 22332
rect 16432 22272 16496 22276
rect 16512 22332 16576 22336
rect 16512 22276 16516 22332
rect 16516 22276 16572 22332
rect 16572 22276 16576 22332
rect 16512 22272 16576 22276
rect 16592 22332 16656 22336
rect 16592 22276 16596 22332
rect 16596 22276 16652 22332
rect 16652 22276 16656 22332
rect 16592 22272 16656 22276
rect 19352 22332 19416 22336
rect 19352 22276 19356 22332
rect 19356 22276 19412 22332
rect 19412 22276 19416 22332
rect 19352 22272 19416 22276
rect 19432 22332 19496 22336
rect 19432 22276 19436 22332
rect 19436 22276 19492 22332
rect 19492 22276 19496 22332
rect 19432 22272 19496 22276
rect 19512 22332 19576 22336
rect 19512 22276 19516 22332
rect 19516 22276 19572 22332
rect 19572 22276 19576 22332
rect 19512 22272 19576 22276
rect 19592 22332 19656 22336
rect 19592 22276 19596 22332
rect 19596 22276 19652 22332
rect 19652 22276 19656 22332
rect 19592 22272 19656 22276
rect 22352 22332 22416 22336
rect 22352 22276 22356 22332
rect 22356 22276 22412 22332
rect 22412 22276 22416 22332
rect 22352 22272 22416 22276
rect 22432 22332 22496 22336
rect 22432 22276 22436 22332
rect 22436 22276 22492 22332
rect 22492 22276 22496 22332
rect 22432 22272 22496 22276
rect 22512 22332 22576 22336
rect 22512 22276 22516 22332
rect 22516 22276 22572 22332
rect 22572 22276 22576 22332
rect 22512 22272 22576 22276
rect 22592 22332 22656 22336
rect 22592 22276 22596 22332
rect 22596 22276 22652 22332
rect 22652 22276 22656 22332
rect 22592 22272 22656 22276
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 2932 21788 2996 21792
rect 2932 21732 2936 21788
rect 2936 21732 2992 21788
rect 2992 21732 2996 21788
rect 2932 21728 2996 21732
rect 3012 21788 3076 21792
rect 3012 21732 3016 21788
rect 3016 21732 3072 21788
rect 3072 21732 3076 21788
rect 3012 21728 3076 21732
rect 3092 21788 3156 21792
rect 3092 21732 3096 21788
rect 3096 21732 3152 21788
rect 3152 21732 3156 21788
rect 3092 21728 3156 21732
rect 5852 21788 5916 21792
rect 5852 21732 5856 21788
rect 5856 21732 5912 21788
rect 5912 21732 5916 21788
rect 5852 21728 5916 21732
rect 5932 21788 5996 21792
rect 5932 21732 5936 21788
rect 5936 21732 5992 21788
rect 5992 21732 5996 21788
rect 5932 21728 5996 21732
rect 6012 21788 6076 21792
rect 6012 21732 6016 21788
rect 6016 21732 6072 21788
rect 6072 21732 6076 21788
rect 6012 21728 6076 21732
rect 6092 21788 6156 21792
rect 6092 21732 6096 21788
rect 6096 21732 6152 21788
rect 6152 21732 6156 21788
rect 6092 21728 6156 21732
rect 8852 21788 8916 21792
rect 8852 21732 8856 21788
rect 8856 21732 8912 21788
rect 8912 21732 8916 21788
rect 8852 21728 8916 21732
rect 8932 21788 8996 21792
rect 8932 21732 8936 21788
rect 8936 21732 8992 21788
rect 8992 21732 8996 21788
rect 8932 21728 8996 21732
rect 9012 21788 9076 21792
rect 9012 21732 9016 21788
rect 9016 21732 9072 21788
rect 9072 21732 9076 21788
rect 9012 21728 9076 21732
rect 9092 21788 9156 21792
rect 9092 21732 9096 21788
rect 9096 21732 9152 21788
rect 9152 21732 9156 21788
rect 9092 21728 9156 21732
rect 11852 21788 11916 21792
rect 11852 21732 11856 21788
rect 11856 21732 11912 21788
rect 11912 21732 11916 21788
rect 11852 21728 11916 21732
rect 11932 21788 11996 21792
rect 11932 21732 11936 21788
rect 11936 21732 11992 21788
rect 11992 21732 11996 21788
rect 11932 21728 11996 21732
rect 12012 21788 12076 21792
rect 12012 21732 12016 21788
rect 12016 21732 12072 21788
rect 12072 21732 12076 21788
rect 12012 21728 12076 21732
rect 12092 21788 12156 21792
rect 12092 21732 12096 21788
rect 12096 21732 12152 21788
rect 12152 21732 12156 21788
rect 12092 21728 12156 21732
rect 14852 21788 14916 21792
rect 14852 21732 14856 21788
rect 14856 21732 14912 21788
rect 14912 21732 14916 21788
rect 14852 21728 14916 21732
rect 14932 21788 14996 21792
rect 14932 21732 14936 21788
rect 14936 21732 14992 21788
rect 14992 21732 14996 21788
rect 14932 21728 14996 21732
rect 15012 21788 15076 21792
rect 15012 21732 15016 21788
rect 15016 21732 15072 21788
rect 15072 21732 15076 21788
rect 15012 21728 15076 21732
rect 15092 21788 15156 21792
rect 15092 21732 15096 21788
rect 15096 21732 15152 21788
rect 15152 21732 15156 21788
rect 15092 21728 15156 21732
rect 17852 21788 17916 21792
rect 17852 21732 17856 21788
rect 17856 21732 17912 21788
rect 17912 21732 17916 21788
rect 17852 21728 17916 21732
rect 17932 21788 17996 21792
rect 17932 21732 17936 21788
rect 17936 21732 17992 21788
rect 17992 21732 17996 21788
rect 17932 21728 17996 21732
rect 18012 21788 18076 21792
rect 18012 21732 18016 21788
rect 18016 21732 18072 21788
rect 18072 21732 18076 21788
rect 18012 21728 18076 21732
rect 18092 21788 18156 21792
rect 18092 21732 18096 21788
rect 18096 21732 18152 21788
rect 18152 21732 18156 21788
rect 18092 21728 18156 21732
rect 20852 21788 20916 21792
rect 20852 21732 20856 21788
rect 20856 21732 20912 21788
rect 20912 21732 20916 21788
rect 20852 21728 20916 21732
rect 20932 21788 20996 21792
rect 20932 21732 20936 21788
rect 20936 21732 20992 21788
rect 20992 21732 20996 21788
rect 20932 21728 20996 21732
rect 21012 21788 21076 21792
rect 21012 21732 21016 21788
rect 21016 21732 21072 21788
rect 21072 21732 21076 21788
rect 21012 21728 21076 21732
rect 21092 21788 21156 21792
rect 21092 21732 21096 21788
rect 21096 21732 21152 21788
rect 21152 21732 21156 21788
rect 21092 21728 21156 21732
rect 23852 21788 23916 21792
rect 23852 21732 23856 21788
rect 23856 21732 23912 21788
rect 23912 21732 23916 21788
rect 23852 21728 23916 21732
rect 23932 21788 23996 21792
rect 23932 21732 23936 21788
rect 23936 21732 23992 21788
rect 23992 21732 23996 21788
rect 23932 21728 23996 21732
rect 24012 21788 24076 21792
rect 24012 21732 24016 21788
rect 24016 21732 24072 21788
rect 24072 21732 24076 21788
rect 24012 21728 24076 21732
rect 24092 21788 24156 21792
rect 24092 21732 24096 21788
rect 24096 21732 24152 21788
rect 24152 21732 24156 21788
rect 24092 21728 24156 21732
rect 1352 21244 1416 21248
rect 1352 21188 1356 21244
rect 1356 21188 1412 21244
rect 1412 21188 1416 21244
rect 1352 21184 1416 21188
rect 1432 21244 1496 21248
rect 1432 21188 1436 21244
rect 1436 21188 1492 21244
rect 1492 21188 1496 21244
rect 1432 21184 1496 21188
rect 1512 21244 1576 21248
rect 1512 21188 1516 21244
rect 1516 21188 1572 21244
rect 1572 21188 1576 21244
rect 1512 21184 1576 21188
rect 1592 21244 1656 21248
rect 1592 21188 1596 21244
rect 1596 21188 1652 21244
rect 1652 21188 1656 21244
rect 1592 21184 1656 21188
rect 4352 21244 4416 21248
rect 4352 21188 4356 21244
rect 4356 21188 4412 21244
rect 4412 21188 4416 21244
rect 4352 21184 4416 21188
rect 4432 21244 4496 21248
rect 4432 21188 4436 21244
rect 4436 21188 4492 21244
rect 4492 21188 4496 21244
rect 4432 21184 4496 21188
rect 4512 21244 4576 21248
rect 4512 21188 4516 21244
rect 4516 21188 4572 21244
rect 4572 21188 4576 21244
rect 4512 21184 4576 21188
rect 4592 21244 4656 21248
rect 4592 21188 4596 21244
rect 4596 21188 4652 21244
rect 4652 21188 4656 21244
rect 4592 21184 4656 21188
rect 7352 21244 7416 21248
rect 7352 21188 7356 21244
rect 7356 21188 7412 21244
rect 7412 21188 7416 21244
rect 7352 21184 7416 21188
rect 7432 21244 7496 21248
rect 7432 21188 7436 21244
rect 7436 21188 7492 21244
rect 7492 21188 7496 21244
rect 7432 21184 7496 21188
rect 7512 21244 7576 21248
rect 7512 21188 7516 21244
rect 7516 21188 7572 21244
rect 7572 21188 7576 21244
rect 7512 21184 7576 21188
rect 7592 21244 7656 21248
rect 7592 21188 7596 21244
rect 7596 21188 7652 21244
rect 7652 21188 7656 21244
rect 7592 21184 7656 21188
rect 10352 21244 10416 21248
rect 10352 21188 10356 21244
rect 10356 21188 10412 21244
rect 10412 21188 10416 21244
rect 10352 21184 10416 21188
rect 10432 21244 10496 21248
rect 10432 21188 10436 21244
rect 10436 21188 10492 21244
rect 10492 21188 10496 21244
rect 10432 21184 10496 21188
rect 10512 21244 10576 21248
rect 10512 21188 10516 21244
rect 10516 21188 10572 21244
rect 10572 21188 10576 21244
rect 10512 21184 10576 21188
rect 10592 21244 10656 21248
rect 10592 21188 10596 21244
rect 10596 21188 10652 21244
rect 10652 21188 10656 21244
rect 10592 21184 10656 21188
rect 13352 21244 13416 21248
rect 13352 21188 13356 21244
rect 13356 21188 13412 21244
rect 13412 21188 13416 21244
rect 13352 21184 13416 21188
rect 13432 21244 13496 21248
rect 13432 21188 13436 21244
rect 13436 21188 13492 21244
rect 13492 21188 13496 21244
rect 13432 21184 13496 21188
rect 13512 21244 13576 21248
rect 13512 21188 13516 21244
rect 13516 21188 13572 21244
rect 13572 21188 13576 21244
rect 13512 21184 13576 21188
rect 13592 21244 13656 21248
rect 13592 21188 13596 21244
rect 13596 21188 13652 21244
rect 13652 21188 13656 21244
rect 13592 21184 13656 21188
rect 16352 21244 16416 21248
rect 16352 21188 16356 21244
rect 16356 21188 16412 21244
rect 16412 21188 16416 21244
rect 16352 21184 16416 21188
rect 16432 21244 16496 21248
rect 16432 21188 16436 21244
rect 16436 21188 16492 21244
rect 16492 21188 16496 21244
rect 16432 21184 16496 21188
rect 16512 21244 16576 21248
rect 16512 21188 16516 21244
rect 16516 21188 16572 21244
rect 16572 21188 16576 21244
rect 16512 21184 16576 21188
rect 16592 21244 16656 21248
rect 16592 21188 16596 21244
rect 16596 21188 16652 21244
rect 16652 21188 16656 21244
rect 16592 21184 16656 21188
rect 19352 21244 19416 21248
rect 19352 21188 19356 21244
rect 19356 21188 19412 21244
rect 19412 21188 19416 21244
rect 19352 21184 19416 21188
rect 19432 21244 19496 21248
rect 19432 21188 19436 21244
rect 19436 21188 19492 21244
rect 19492 21188 19496 21244
rect 19432 21184 19496 21188
rect 19512 21244 19576 21248
rect 19512 21188 19516 21244
rect 19516 21188 19572 21244
rect 19572 21188 19576 21244
rect 19512 21184 19576 21188
rect 19592 21244 19656 21248
rect 19592 21188 19596 21244
rect 19596 21188 19652 21244
rect 19652 21188 19656 21244
rect 19592 21184 19656 21188
rect 22352 21244 22416 21248
rect 22352 21188 22356 21244
rect 22356 21188 22412 21244
rect 22412 21188 22416 21244
rect 22352 21184 22416 21188
rect 22432 21244 22496 21248
rect 22432 21188 22436 21244
rect 22436 21188 22492 21244
rect 22492 21188 22496 21244
rect 22432 21184 22496 21188
rect 22512 21244 22576 21248
rect 22512 21188 22516 21244
rect 22516 21188 22572 21244
rect 22572 21188 22576 21244
rect 22512 21184 22576 21188
rect 22592 21244 22656 21248
rect 22592 21188 22596 21244
rect 22596 21188 22652 21244
rect 22652 21188 22656 21244
rect 22592 21184 22656 21188
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 2932 20700 2996 20704
rect 2932 20644 2936 20700
rect 2936 20644 2992 20700
rect 2992 20644 2996 20700
rect 2932 20640 2996 20644
rect 3012 20700 3076 20704
rect 3012 20644 3016 20700
rect 3016 20644 3072 20700
rect 3072 20644 3076 20700
rect 3012 20640 3076 20644
rect 3092 20700 3156 20704
rect 3092 20644 3096 20700
rect 3096 20644 3152 20700
rect 3152 20644 3156 20700
rect 3092 20640 3156 20644
rect 5852 20700 5916 20704
rect 5852 20644 5856 20700
rect 5856 20644 5912 20700
rect 5912 20644 5916 20700
rect 5852 20640 5916 20644
rect 5932 20700 5996 20704
rect 5932 20644 5936 20700
rect 5936 20644 5992 20700
rect 5992 20644 5996 20700
rect 5932 20640 5996 20644
rect 6012 20700 6076 20704
rect 6012 20644 6016 20700
rect 6016 20644 6072 20700
rect 6072 20644 6076 20700
rect 6012 20640 6076 20644
rect 6092 20700 6156 20704
rect 6092 20644 6096 20700
rect 6096 20644 6152 20700
rect 6152 20644 6156 20700
rect 6092 20640 6156 20644
rect 8852 20700 8916 20704
rect 8852 20644 8856 20700
rect 8856 20644 8912 20700
rect 8912 20644 8916 20700
rect 8852 20640 8916 20644
rect 8932 20700 8996 20704
rect 8932 20644 8936 20700
rect 8936 20644 8992 20700
rect 8992 20644 8996 20700
rect 8932 20640 8996 20644
rect 9012 20700 9076 20704
rect 9012 20644 9016 20700
rect 9016 20644 9072 20700
rect 9072 20644 9076 20700
rect 9012 20640 9076 20644
rect 9092 20700 9156 20704
rect 9092 20644 9096 20700
rect 9096 20644 9152 20700
rect 9152 20644 9156 20700
rect 9092 20640 9156 20644
rect 11852 20700 11916 20704
rect 11852 20644 11856 20700
rect 11856 20644 11912 20700
rect 11912 20644 11916 20700
rect 11852 20640 11916 20644
rect 11932 20700 11996 20704
rect 11932 20644 11936 20700
rect 11936 20644 11992 20700
rect 11992 20644 11996 20700
rect 11932 20640 11996 20644
rect 12012 20700 12076 20704
rect 12012 20644 12016 20700
rect 12016 20644 12072 20700
rect 12072 20644 12076 20700
rect 12012 20640 12076 20644
rect 12092 20700 12156 20704
rect 12092 20644 12096 20700
rect 12096 20644 12152 20700
rect 12152 20644 12156 20700
rect 12092 20640 12156 20644
rect 14852 20700 14916 20704
rect 14852 20644 14856 20700
rect 14856 20644 14912 20700
rect 14912 20644 14916 20700
rect 14852 20640 14916 20644
rect 14932 20700 14996 20704
rect 14932 20644 14936 20700
rect 14936 20644 14992 20700
rect 14992 20644 14996 20700
rect 14932 20640 14996 20644
rect 15012 20700 15076 20704
rect 15012 20644 15016 20700
rect 15016 20644 15072 20700
rect 15072 20644 15076 20700
rect 15012 20640 15076 20644
rect 15092 20700 15156 20704
rect 15092 20644 15096 20700
rect 15096 20644 15152 20700
rect 15152 20644 15156 20700
rect 15092 20640 15156 20644
rect 17852 20700 17916 20704
rect 17852 20644 17856 20700
rect 17856 20644 17912 20700
rect 17912 20644 17916 20700
rect 17852 20640 17916 20644
rect 17932 20700 17996 20704
rect 17932 20644 17936 20700
rect 17936 20644 17992 20700
rect 17992 20644 17996 20700
rect 17932 20640 17996 20644
rect 18012 20700 18076 20704
rect 18012 20644 18016 20700
rect 18016 20644 18072 20700
rect 18072 20644 18076 20700
rect 18012 20640 18076 20644
rect 18092 20700 18156 20704
rect 18092 20644 18096 20700
rect 18096 20644 18152 20700
rect 18152 20644 18156 20700
rect 18092 20640 18156 20644
rect 20852 20700 20916 20704
rect 20852 20644 20856 20700
rect 20856 20644 20912 20700
rect 20912 20644 20916 20700
rect 20852 20640 20916 20644
rect 20932 20700 20996 20704
rect 20932 20644 20936 20700
rect 20936 20644 20992 20700
rect 20992 20644 20996 20700
rect 20932 20640 20996 20644
rect 21012 20700 21076 20704
rect 21012 20644 21016 20700
rect 21016 20644 21072 20700
rect 21072 20644 21076 20700
rect 21012 20640 21076 20644
rect 21092 20700 21156 20704
rect 21092 20644 21096 20700
rect 21096 20644 21152 20700
rect 21152 20644 21156 20700
rect 21092 20640 21156 20644
rect 23852 20700 23916 20704
rect 23852 20644 23856 20700
rect 23856 20644 23912 20700
rect 23912 20644 23916 20700
rect 23852 20640 23916 20644
rect 23932 20700 23996 20704
rect 23932 20644 23936 20700
rect 23936 20644 23992 20700
rect 23992 20644 23996 20700
rect 23932 20640 23996 20644
rect 24012 20700 24076 20704
rect 24012 20644 24016 20700
rect 24016 20644 24072 20700
rect 24072 20644 24076 20700
rect 24012 20640 24076 20644
rect 24092 20700 24156 20704
rect 24092 20644 24096 20700
rect 24096 20644 24152 20700
rect 24152 20644 24156 20700
rect 24092 20640 24156 20644
rect 1352 20156 1416 20160
rect 1352 20100 1356 20156
rect 1356 20100 1412 20156
rect 1412 20100 1416 20156
rect 1352 20096 1416 20100
rect 1432 20156 1496 20160
rect 1432 20100 1436 20156
rect 1436 20100 1492 20156
rect 1492 20100 1496 20156
rect 1432 20096 1496 20100
rect 1512 20156 1576 20160
rect 1512 20100 1516 20156
rect 1516 20100 1572 20156
rect 1572 20100 1576 20156
rect 1512 20096 1576 20100
rect 1592 20156 1656 20160
rect 1592 20100 1596 20156
rect 1596 20100 1652 20156
rect 1652 20100 1656 20156
rect 1592 20096 1656 20100
rect 4352 20156 4416 20160
rect 4352 20100 4356 20156
rect 4356 20100 4412 20156
rect 4412 20100 4416 20156
rect 4352 20096 4416 20100
rect 4432 20156 4496 20160
rect 4432 20100 4436 20156
rect 4436 20100 4492 20156
rect 4492 20100 4496 20156
rect 4432 20096 4496 20100
rect 4512 20156 4576 20160
rect 4512 20100 4516 20156
rect 4516 20100 4572 20156
rect 4572 20100 4576 20156
rect 4512 20096 4576 20100
rect 4592 20156 4656 20160
rect 4592 20100 4596 20156
rect 4596 20100 4652 20156
rect 4652 20100 4656 20156
rect 4592 20096 4656 20100
rect 7352 20156 7416 20160
rect 7352 20100 7356 20156
rect 7356 20100 7412 20156
rect 7412 20100 7416 20156
rect 7352 20096 7416 20100
rect 7432 20156 7496 20160
rect 7432 20100 7436 20156
rect 7436 20100 7492 20156
rect 7492 20100 7496 20156
rect 7432 20096 7496 20100
rect 7512 20156 7576 20160
rect 7512 20100 7516 20156
rect 7516 20100 7572 20156
rect 7572 20100 7576 20156
rect 7512 20096 7576 20100
rect 7592 20156 7656 20160
rect 7592 20100 7596 20156
rect 7596 20100 7652 20156
rect 7652 20100 7656 20156
rect 7592 20096 7656 20100
rect 10352 20156 10416 20160
rect 10352 20100 10356 20156
rect 10356 20100 10412 20156
rect 10412 20100 10416 20156
rect 10352 20096 10416 20100
rect 10432 20156 10496 20160
rect 10432 20100 10436 20156
rect 10436 20100 10492 20156
rect 10492 20100 10496 20156
rect 10432 20096 10496 20100
rect 10512 20156 10576 20160
rect 10512 20100 10516 20156
rect 10516 20100 10572 20156
rect 10572 20100 10576 20156
rect 10512 20096 10576 20100
rect 10592 20156 10656 20160
rect 10592 20100 10596 20156
rect 10596 20100 10652 20156
rect 10652 20100 10656 20156
rect 10592 20096 10656 20100
rect 13352 20156 13416 20160
rect 13352 20100 13356 20156
rect 13356 20100 13412 20156
rect 13412 20100 13416 20156
rect 13352 20096 13416 20100
rect 13432 20156 13496 20160
rect 13432 20100 13436 20156
rect 13436 20100 13492 20156
rect 13492 20100 13496 20156
rect 13432 20096 13496 20100
rect 13512 20156 13576 20160
rect 13512 20100 13516 20156
rect 13516 20100 13572 20156
rect 13572 20100 13576 20156
rect 13512 20096 13576 20100
rect 13592 20156 13656 20160
rect 13592 20100 13596 20156
rect 13596 20100 13652 20156
rect 13652 20100 13656 20156
rect 13592 20096 13656 20100
rect 16352 20156 16416 20160
rect 16352 20100 16356 20156
rect 16356 20100 16412 20156
rect 16412 20100 16416 20156
rect 16352 20096 16416 20100
rect 16432 20156 16496 20160
rect 16432 20100 16436 20156
rect 16436 20100 16492 20156
rect 16492 20100 16496 20156
rect 16432 20096 16496 20100
rect 16512 20156 16576 20160
rect 16512 20100 16516 20156
rect 16516 20100 16572 20156
rect 16572 20100 16576 20156
rect 16512 20096 16576 20100
rect 16592 20156 16656 20160
rect 16592 20100 16596 20156
rect 16596 20100 16652 20156
rect 16652 20100 16656 20156
rect 16592 20096 16656 20100
rect 19352 20156 19416 20160
rect 19352 20100 19356 20156
rect 19356 20100 19412 20156
rect 19412 20100 19416 20156
rect 19352 20096 19416 20100
rect 19432 20156 19496 20160
rect 19432 20100 19436 20156
rect 19436 20100 19492 20156
rect 19492 20100 19496 20156
rect 19432 20096 19496 20100
rect 19512 20156 19576 20160
rect 19512 20100 19516 20156
rect 19516 20100 19572 20156
rect 19572 20100 19576 20156
rect 19512 20096 19576 20100
rect 19592 20156 19656 20160
rect 19592 20100 19596 20156
rect 19596 20100 19652 20156
rect 19652 20100 19656 20156
rect 19592 20096 19656 20100
rect 22352 20156 22416 20160
rect 22352 20100 22356 20156
rect 22356 20100 22412 20156
rect 22412 20100 22416 20156
rect 22352 20096 22416 20100
rect 22432 20156 22496 20160
rect 22432 20100 22436 20156
rect 22436 20100 22492 20156
rect 22492 20100 22496 20156
rect 22432 20096 22496 20100
rect 22512 20156 22576 20160
rect 22512 20100 22516 20156
rect 22516 20100 22572 20156
rect 22572 20100 22576 20156
rect 22512 20096 22576 20100
rect 22592 20156 22656 20160
rect 22592 20100 22596 20156
rect 22596 20100 22652 20156
rect 22652 20100 22656 20156
rect 22592 20096 22656 20100
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 2932 19612 2996 19616
rect 2932 19556 2936 19612
rect 2936 19556 2992 19612
rect 2992 19556 2996 19612
rect 2932 19552 2996 19556
rect 3012 19612 3076 19616
rect 3012 19556 3016 19612
rect 3016 19556 3072 19612
rect 3072 19556 3076 19612
rect 3012 19552 3076 19556
rect 3092 19612 3156 19616
rect 3092 19556 3096 19612
rect 3096 19556 3152 19612
rect 3152 19556 3156 19612
rect 3092 19552 3156 19556
rect 5852 19612 5916 19616
rect 5852 19556 5856 19612
rect 5856 19556 5912 19612
rect 5912 19556 5916 19612
rect 5852 19552 5916 19556
rect 5932 19612 5996 19616
rect 5932 19556 5936 19612
rect 5936 19556 5992 19612
rect 5992 19556 5996 19612
rect 5932 19552 5996 19556
rect 6012 19612 6076 19616
rect 6012 19556 6016 19612
rect 6016 19556 6072 19612
rect 6072 19556 6076 19612
rect 6012 19552 6076 19556
rect 6092 19612 6156 19616
rect 6092 19556 6096 19612
rect 6096 19556 6152 19612
rect 6152 19556 6156 19612
rect 6092 19552 6156 19556
rect 8852 19612 8916 19616
rect 8852 19556 8856 19612
rect 8856 19556 8912 19612
rect 8912 19556 8916 19612
rect 8852 19552 8916 19556
rect 8932 19612 8996 19616
rect 8932 19556 8936 19612
rect 8936 19556 8992 19612
rect 8992 19556 8996 19612
rect 8932 19552 8996 19556
rect 9012 19612 9076 19616
rect 9012 19556 9016 19612
rect 9016 19556 9072 19612
rect 9072 19556 9076 19612
rect 9012 19552 9076 19556
rect 9092 19612 9156 19616
rect 9092 19556 9096 19612
rect 9096 19556 9152 19612
rect 9152 19556 9156 19612
rect 9092 19552 9156 19556
rect 11852 19612 11916 19616
rect 11852 19556 11856 19612
rect 11856 19556 11912 19612
rect 11912 19556 11916 19612
rect 11852 19552 11916 19556
rect 11932 19612 11996 19616
rect 11932 19556 11936 19612
rect 11936 19556 11992 19612
rect 11992 19556 11996 19612
rect 11932 19552 11996 19556
rect 12012 19612 12076 19616
rect 12012 19556 12016 19612
rect 12016 19556 12072 19612
rect 12072 19556 12076 19612
rect 12012 19552 12076 19556
rect 12092 19612 12156 19616
rect 12092 19556 12096 19612
rect 12096 19556 12152 19612
rect 12152 19556 12156 19612
rect 12092 19552 12156 19556
rect 14852 19612 14916 19616
rect 14852 19556 14856 19612
rect 14856 19556 14912 19612
rect 14912 19556 14916 19612
rect 14852 19552 14916 19556
rect 14932 19612 14996 19616
rect 14932 19556 14936 19612
rect 14936 19556 14992 19612
rect 14992 19556 14996 19612
rect 14932 19552 14996 19556
rect 15012 19612 15076 19616
rect 15012 19556 15016 19612
rect 15016 19556 15072 19612
rect 15072 19556 15076 19612
rect 15012 19552 15076 19556
rect 15092 19612 15156 19616
rect 15092 19556 15096 19612
rect 15096 19556 15152 19612
rect 15152 19556 15156 19612
rect 15092 19552 15156 19556
rect 17852 19612 17916 19616
rect 17852 19556 17856 19612
rect 17856 19556 17912 19612
rect 17912 19556 17916 19612
rect 17852 19552 17916 19556
rect 17932 19612 17996 19616
rect 17932 19556 17936 19612
rect 17936 19556 17992 19612
rect 17992 19556 17996 19612
rect 17932 19552 17996 19556
rect 18012 19612 18076 19616
rect 18012 19556 18016 19612
rect 18016 19556 18072 19612
rect 18072 19556 18076 19612
rect 18012 19552 18076 19556
rect 18092 19612 18156 19616
rect 18092 19556 18096 19612
rect 18096 19556 18152 19612
rect 18152 19556 18156 19612
rect 18092 19552 18156 19556
rect 20852 19612 20916 19616
rect 20852 19556 20856 19612
rect 20856 19556 20912 19612
rect 20912 19556 20916 19612
rect 20852 19552 20916 19556
rect 20932 19612 20996 19616
rect 20932 19556 20936 19612
rect 20936 19556 20992 19612
rect 20992 19556 20996 19612
rect 20932 19552 20996 19556
rect 21012 19612 21076 19616
rect 21012 19556 21016 19612
rect 21016 19556 21072 19612
rect 21072 19556 21076 19612
rect 21012 19552 21076 19556
rect 21092 19612 21156 19616
rect 21092 19556 21096 19612
rect 21096 19556 21152 19612
rect 21152 19556 21156 19612
rect 21092 19552 21156 19556
rect 23852 19612 23916 19616
rect 23852 19556 23856 19612
rect 23856 19556 23912 19612
rect 23912 19556 23916 19612
rect 23852 19552 23916 19556
rect 23932 19612 23996 19616
rect 23932 19556 23936 19612
rect 23936 19556 23992 19612
rect 23992 19556 23996 19612
rect 23932 19552 23996 19556
rect 24012 19612 24076 19616
rect 24012 19556 24016 19612
rect 24016 19556 24072 19612
rect 24072 19556 24076 19612
rect 24012 19552 24076 19556
rect 24092 19612 24156 19616
rect 24092 19556 24096 19612
rect 24096 19556 24152 19612
rect 24152 19556 24156 19612
rect 24092 19552 24156 19556
rect 1352 19068 1416 19072
rect 1352 19012 1356 19068
rect 1356 19012 1412 19068
rect 1412 19012 1416 19068
rect 1352 19008 1416 19012
rect 1432 19068 1496 19072
rect 1432 19012 1436 19068
rect 1436 19012 1492 19068
rect 1492 19012 1496 19068
rect 1432 19008 1496 19012
rect 1512 19068 1576 19072
rect 1512 19012 1516 19068
rect 1516 19012 1572 19068
rect 1572 19012 1576 19068
rect 1512 19008 1576 19012
rect 1592 19068 1656 19072
rect 1592 19012 1596 19068
rect 1596 19012 1652 19068
rect 1652 19012 1656 19068
rect 1592 19008 1656 19012
rect 4352 19068 4416 19072
rect 4352 19012 4356 19068
rect 4356 19012 4412 19068
rect 4412 19012 4416 19068
rect 4352 19008 4416 19012
rect 4432 19068 4496 19072
rect 4432 19012 4436 19068
rect 4436 19012 4492 19068
rect 4492 19012 4496 19068
rect 4432 19008 4496 19012
rect 4512 19068 4576 19072
rect 4512 19012 4516 19068
rect 4516 19012 4572 19068
rect 4572 19012 4576 19068
rect 4512 19008 4576 19012
rect 4592 19068 4656 19072
rect 4592 19012 4596 19068
rect 4596 19012 4652 19068
rect 4652 19012 4656 19068
rect 4592 19008 4656 19012
rect 7352 19068 7416 19072
rect 7352 19012 7356 19068
rect 7356 19012 7412 19068
rect 7412 19012 7416 19068
rect 7352 19008 7416 19012
rect 7432 19068 7496 19072
rect 7432 19012 7436 19068
rect 7436 19012 7492 19068
rect 7492 19012 7496 19068
rect 7432 19008 7496 19012
rect 7512 19068 7576 19072
rect 7512 19012 7516 19068
rect 7516 19012 7572 19068
rect 7572 19012 7576 19068
rect 7512 19008 7576 19012
rect 7592 19068 7656 19072
rect 7592 19012 7596 19068
rect 7596 19012 7652 19068
rect 7652 19012 7656 19068
rect 7592 19008 7656 19012
rect 10352 19068 10416 19072
rect 10352 19012 10356 19068
rect 10356 19012 10412 19068
rect 10412 19012 10416 19068
rect 10352 19008 10416 19012
rect 10432 19068 10496 19072
rect 10432 19012 10436 19068
rect 10436 19012 10492 19068
rect 10492 19012 10496 19068
rect 10432 19008 10496 19012
rect 10512 19068 10576 19072
rect 10512 19012 10516 19068
rect 10516 19012 10572 19068
rect 10572 19012 10576 19068
rect 10512 19008 10576 19012
rect 10592 19068 10656 19072
rect 10592 19012 10596 19068
rect 10596 19012 10652 19068
rect 10652 19012 10656 19068
rect 10592 19008 10656 19012
rect 13352 19068 13416 19072
rect 13352 19012 13356 19068
rect 13356 19012 13412 19068
rect 13412 19012 13416 19068
rect 13352 19008 13416 19012
rect 13432 19068 13496 19072
rect 13432 19012 13436 19068
rect 13436 19012 13492 19068
rect 13492 19012 13496 19068
rect 13432 19008 13496 19012
rect 13512 19068 13576 19072
rect 13512 19012 13516 19068
rect 13516 19012 13572 19068
rect 13572 19012 13576 19068
rect 13512 19008 13576 19012
rect 13592 19068 13656 19072
rect 13592 19012 13596 19068
rect 13596 19012 13652 19068
rect 13652 19012 13656 19068
rect 13592 19008 13656 19012
rect 16352 19068 16416 19072
rect 16352 19012 16356 19068
rect 16356 19012 16412 19068
rect 16412 19012 16416 19068
rect 16352 19008 16416 19012
rect 16432 19068 16496 19072
rect 16432 19012 16436 19068
rect 16436 19012 16492 19068
rect 16492 19012 16496 19068
rect 16432 19008 16496 19012
rect 16512 19068 16576 19072
rect 16512 19012 16516 19068
rect 16516 19012 16572 19068
rect 16572 19012 16576 19068
rect 16512 19008 16576 19012
rect 16592 19068 16656 19072
rect 16592 19012 16596 19068
rect 16596 19012 16652 19068
rect 16652 19012 16656 19068
rect 16592 19008 16656 19012
rect 19352 19068 19416 19072
rect 19352 19012 19356 19068
rect 19356 19012 19412 19068
rect 19412 19012 19416 19068
rect 19352 19008 19416 19012
rect 19432 19068 19496 19072
rect 19432 19012 19436 19068
rect 19436 19012 19492 19068
rect 19492 19012 19496 19068
rect 19432 19008 19496 19012
rect 19512 19068 19576 19072
rect 19512 19012 19516 19068
rect 19516 19012 19572 19068
rect 19572 19012 19576 19068
rect 19512 19008 19576 19012
rect 19592 19068 19656 19072
rect 19592 19012 19596 19068
rect 19596 19012 19652 19068
rect 19652 19012 19656 19068
rect 19592 19008 19656 19012
rect 22352 19068 22416 19072
rect 22352 19012 22356 19068
rect 22356 19012 22412 19068
rect 22412 19012 22416 19068
rect 22352 19008 22416 19012
rect 22432 19068 22496 19072
rect 22432 19012 22436 19068
rect 22436 19012 22492 19068
rect 22492 19012 22496 19068
rect 22432 19008 22496 19012
rect 22512 19068 22576 19072
rect 22512 19012 22516 19068
rect 22516 19012 22572 19068
rect 22572 19012 22576 19068
rect 22512 19008 22576 19012
rect 22592 19068 22656 19072
rect 22592 19012 22596 19068
rect 22596 19012 22652 19068
rect 22652 19012 22656 19068
rect 22592 19008 22656 19012
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 2932 18524 2996 18528
rect 2932 18468 2936 18524
rect 2936 18468 2992 18524
rect 2992 18468 2996 18524
rect 2932 18464 2996 18468
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 5852 18524 5916 18528
rect 5852 18468 5856 18524
rect 5856 18468 5912 18524
rect 5912 18468 5916 18524
rect 5852 18464 5916 18468
rect 5932 18524 5996 18528
rect 5932 18468 5936 18524
rect 5936 18468 5992 18524
rect 5992 18468 5996 18524
rect 5932 18464 5996 18468
rect 6012 18524 6076 18528
rect 6012 18468 6016 18524
rect 6016 18468 6072 18524
rect 6072 18468 6076 18524
rect 6012 18464 6076 18468
rect 6092 18524 6156 18528
rect 6092 18468 6096 18524
rect 6096 18468 6152 18524
rect 6152 18468 6156 18524
rect 6092 18464 6156 18468
rect 8852 18524 8916 18528
rect 8852 18468 8856 18524
rect 8856 18468 8912 18524
rect 8912 18468 8916 18524
rect 8852 18464 8916 18468
rect 8932 18524 8996 18528
rect 8932 18468 8936 18524
rect 8936 18468 8992 18524
rect 8992 18468 8996 18524
rect 8932 18464 8996 18468
rect 9012 18524 9076 18528
rect 9012 18468 9016 18524
rect 9016 18468 9072 18524
rect 9072 18468 9076 18524
rect 9012 18464 9076 18468
rect 9092 18524 9156 18528
rect 9092 18468 9096 18524
rect 9096 18468 9152 18524
rect 9152 18468 9156 18524
rect 9092 18464 9156 18468
rect 11852 18524 11916 18528
rect 11852 18468 11856 18524
rect 11856 18468 11912 18524
rect 11912 18468 11916 18524
rect 11852 18464 11916 18468
rect 11932 18524 11996 18528
rect 11932 18468 11936 18524
rect 11936 18468 11992 18524
rect 11992 18468 11996 18524
rect 11932 18464 11996 18468
rect 12012 18524 12076 18528
rect 12012 18468 12016 18524
rect 12016 18468 12072 18524
rect 12072 18468 12076 18524
rect 12012 18464 12076 18468
rect 12092 18524 12156 18528
rect 12092 18468 12096 18524
rect 12096 18468 12152 18524
rect 12152 18468 12156 18524
rect 12092 18464 12156 18468
rect 14852 18524 14916 18528
rect 14852 18468 14856 18524
rect 14856 18468 14912 18524
rect 14912 18468 14916 18524
rect 14852 18464 14916 18468
rect 14932 18524 14996 18528
rect 14932 18468 14936 18524
rect 14936 18468 14992 18524
rect 14992 18468 14996 18524
rect 14932 18464 14996 18468
rect 15012 18524 15076 18528
rect 15012 18468 15016 18524
rect 15016 18468 15072 18524
rect 15072 18468 15076 18524
rect 15012 18464 15076 18468
rect 15092 18524 15156 18528
rect 15092 18468 15096 18524
rect 15096 18468 15152 18524
rect 15152 18468 15156 18524
rect 15092 18464 15156 18468
rect 17852 18524 17916 18528
rect 17852 18468 17856 18524
rect 17856 18468 17912 18524
rect 17912 18468 17916 18524
rect 17852 18464 17916 18468
rect 17932 18524 17996 18528
rect 17932 18468 17936 18524
rect 17936 18468 17992 18524
rect 17992 18468 17996 18524
rect 17932 18464 17996 18468
rect 18012 18524 18076 18528
rect 18012 18468 18016 18524
rect 18016 18468 18072 18524
rect 18072 18468 18076 18524
rect 18012 18464 18076 18468
rect 18092 18524 18156 18528
rect 18092 18468 18096 18524
rect 18096 18468 18152 18524
rect 18152 18468 18156 18524
rect 18092 18464 18156 18468
rect 20852 18524 20916 18528
rect 20852 18468 20856 18524
rect 20856 18468 20912 18524
rect 20912 18468 20916 18524
rect 20852 18464 20916 18468
rect 20932 18524 20996 18528
rect 20932 18468 20936 18524
rect 20936 18468 20992 18524
rect 20992 18468 20996 18524
rect 20932 18464 20996 18468
rect 21012 18524 21076 18528
rect 21012 18468 21016 18524
rect 21016 18468 21072 18524
rect 21072 18468 21076 18524
rect 21012 18464 21076 18468
rect 21092 18524 21156 18528
rect 21092 18468 21096 18524
rect 21096 18468 21152 18524
rect 21152 18468 21156 18524
rect 21092 18464 21156 18468
rect 23852 18524 23916 18528
rect 23852 18468 23856 18524
rect 23856 18468 23912 18524
rect 23912 18468 23916 18524
rect 23852 18464 23916 18468
rect 23932 18524 23996 18528
rect 23932 18468 23936 18524
rect 23936 18468 23992 18524
rect 23992 18468 23996 18524
rect 23932 18464 23996 18468
rect 24012 18524 24076 18528
rect 24012 18468 24016 18524
rect 24016 18468 24072 18524
rect 24072 18468 24076 18524
rect 24012 18464 24076 18468
rect 24092 18524 24156 18528
rect 24092 18468 24096 18524
rect 24096 18468 24152 18524
rect 24152 18468 24156 18524
rect 24092 18464 24156 18468
rect 13124 18260 13188 18324
rect 1352 17980 1416 17984
rect 1352 17924 1356 17980
rect 1356 17924 1412 17980
rect 1412 17924 1416 17980
rect 1352 17920 1416 17924
rect 1432 17980 1496 17984
rect 1432 17924 1436 17980
rect 1436 17924 1492 17980
rect 1492 17924 1496 17980
rect 1432 17920 1496 17924
rect 1512 17980 1576 17984
rect 1512 17924 1516 17980
rect 1516 17924 1572 17980
rect 1572 17924 1576 17980
rect 1512 17920 1576 17924
rect 1592 17980 1656 17984
rect 1592 17924 1596 17980
rect 1596 17924 1652 17980
rect 1652 17924 1656 17980
rect 1592 17920 1656 17924
rect 4352 17980 4416 17984
rect 4352 17924 4356 17980
rect 4356 17924 4412 17980
rect 4412 17924 4416 17980
rect 4352 17920 4416 17924
rect 4432 17980 4496 17984
rect 4432 17924 4436 17980
rect 4436 17924 4492 17980
rect 4492 17924 4496 17980
rect 4432 17920 4496 17924
rect 4512 17980 4576 17984
rect 4512 17924 4516 17980
rect 4516 17924 4572 17980
rect 4572 17924 4576 17980
rect 4512 17920 4576 17924
rect 4592 17980 4656 17984
rect 4592 17924 4596 17980
rect 4596 17924 4652 17980
rect 4652 17924 4656 17980
rect 4592 17920 4656 17924
rect 7352 17980 7416 17984
rect 7352 17924 7356 17980
rect 7356 17924 7412 17980
rect 7412 17924 7416 17980
rect 7352 17920 7416 17924
rect 7432 17980 7496 17984
rect 7432 17924 7436 17980
rect 7436 17924 7492 17980
rect 7492 17924 7496 17980
rect 7432 17920 7496 17924
rect 7512 17980 7576 17984
rect 7512 17924 7516 17980
rect 7516 17924 7572 17980
rect 7572 17924 7576 17980
rect 7512 17920 7576 17924
rect 7592 17980 7656 17984
rect 7592 17924 7596 17980
rect 7596 17924 7652 17980
rect 7652 17924 7656 17980
rect 7592 17920 7656 17924
rect 10352 17980 10416 17984
rect 10352 17924 10356 17980
rect 10356 17924 10412 17980
rect 10412 17924 10416 17980
rect 10352 17920 10416 17924
rect 10432 17980 10496 17984
rect 10432 17924 10436 17980
rect 10436 17924 10492 17980
rect 10492 17924 10496 17980
rect 10432 17920 10496 17924
rect 10512 17980 10576 17984
rect 10512 17924 10516 17980
rect 10516 17924 10572 17980
rect 10572 17924 10576 17980
rect 10512 17920 10576 17924
rect 10592 17980 10656 17984
rect 10592 17924 10596 17980
rect 10596 17924 10652 17980
rect 10652 17924 10656 17980
rect 10592 17920 10656 17924
rect 13352 17980 13416 17984
rect 13352 17924 13356 17980
rect 13356 17924 13412 17980
rect 13412 17924 13416 17980
rect 13352 17920 13416 17924
rect 13432 17980 13496 17984
rect 13432 17924 13436 17980
rect 13436 17924 13492 17980
rect 13492 17924 13496 17980
rect 13432 17920 13496 17924
rect 13512 17980 13576 17984
rect 13512 17924 13516 17980
rect 13516 17924 13572 17980
rect 13572 17924 13576 17980
rect 13512 17920 13576 17924
rect 13592 17980 13656 17984
rect 13592 17924 13596 17980
rect 13596 17924 13652 17980
rect 13652 17924 13656 17980
rect 13592 17920 13656 17924
rect 16352 17980 16416 17984
rect 16352 17924 16356 17980
rect 16356 17924 16412 17980
rect 16412 17924 16416 17980
rect 16352 17920 16416 17924
rect 16432 17980 16496 17984
rect 16432 17924 16436 17980
rect 16436 17924 16492 17980
rect 16492 17924 16496 17980
rect 16432 17920 16496 17924
rect 16512 17980 16576 17984
rect 16512 17924 16516 17980
rect 16516 17924 16572 17980
rect 16572 17924 16576 17980
rect 16512 17920 16576 17924
rect 16592 17980 16656 17984
rect 16592 17924 16596 17980
rect 16596 17924 16652 17980
rect 16652 17924 16656 17980
rect 16592 17920 16656 17924
rect 19352 17980 19416 17984
rect 19352 17924 19356 17980
rect 19356 17924 19412 17980
rect 19412 17924 19416 17980
rect 19352 17920 19416 17924
rect 19432 17980 19496 17984
rect 19432 17924 19436 17980
rect 19436 17924 19492 17980
rect 19492 17924 19496 17980
rect 19432 17920 19496 17924
rect 19512 17980 19576 17984
rect 19512 17924 19516 17980
rect 19516 17924 19572 17980
rect 19572 17924 19576 17980
rect 19512 17920 19576 17924
rect 19592 17980 19656 17984
rect 19592 17924 19596 17980
rect 19596 17924 19652 17980
rect 19652 17924 19656 17980
rect 19592 17920 19656 17924
rect 22140 18124 22204 18188
rect 22352 17980 22416 17984
rect 22352 17924 22356 17980
rect 22356 17924 22412 17980
rect 22412 17924 22416 17980
rect 22352 17920 22416 17924
rect 22432 17980 22496 17984
rect 22432 17924 22436 17980
rect 22436 17924 22492 17980
rect 22492 17924 22496 17980
rect 22432 17920 22496 17924
rect 22512 17980 22576 17984
rect 22512 17924 22516 17980
rect 22516 17924 22572 17980
rect 22572 17924 22576 17980
rect 22512 17920 22576 17924
rect 22592 17980 22656 17984
rect 22592 17924 22596 17980
rect 22596 17924 22652 17980
rect 22652 17924 22656 17980
rect 22592 17920 22656 17924
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 2932 17436 2996 17440
rect 2932 17380 2936 17436
rect 2936 17380 2992 17436
rect 2992 17380 2996 17436
rect 2932 17376 2996 17380
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 5852 17436 5916 17440
rect 5852 17380 5856 17436
rect 5856 17380 5912 17436
rect 5912 17380 5916 17436
rect 5852 17376 5916 17380
rect 5932 17436 5996 17440
rect 5932 17380 5936 17436
rect 5936 17380 5992 17436
rect 5992 17380 5996 17436
rect 5932 17376 5996 17380
rect 6012 17436 6076 17440
rect 6012 17380 6016 17436
rect 6016 17380 6072 17436
rect 6072 17380 6076 17436
rect 6012 17376 6076 17380
rect 6092 17436 6156 17440
rect 6092 17380 6096 17436
rect 6096 17380 6152 17436
rect 6152 17380 6156 17436
rect 6092 17376 6156 17380
rect 8852 17436 8916 17440
rect 8852 17380 8856 17436
rect 8856 17380 8912 17436
rect 8912 17380 8916 17436
rect 8852 17376 8916 17380
rect 8932 17436 8996 17440
rect 8932 17380 8936 17436
rect 8936 17380 8992 17436
rect 8992 17380 8996 17436
rect 8932 17376 8996 17380
rect 9012 17436 9076 17440
rect 9012 17380 9016 17436
rect 9016 17380 9072 17436
rect 9072 17380 9076 17436
rect 9012 17376 9076 17380
rect 9092 17436 9156 17440
rect 9092 17380 9096 17436
rect 9096 17380 9152 17436
rect 9152 17380 9156 17436
rect 9092 17376 9156 17380
rect 11852 17436 11916 17440
rect 11852 17380 11856 17436
rect 11856 17380 11912 17436
rect 11912 17380 11916 17436
rect 11852 17376 11916 17380
rect 11932 17436 11996 17440
rect 11932 17380 11936 17436
rect 11936 17380 11992 17436
rect 11992 17380 11996 17436
rect 11932 17376 11996 17380
rect 12012 17436 12076 17440
rect 12012 17380 12016 17436
rect 12016 17380 12072 17436
rect 12072 17380 12076 17436
rect 12012 17376 12076 17380
rect 12092 17436 12156 17440
rect 12092 17380 12096 17436
rect 12096 17380 12152 17436
rect 12152 17380 12156 17436
rect 12092 17376 12156 17380
rect 14852 17436 14916 17440
rect 14852 17380 14856 17436
rect 14856 17380 14912 17436
rect 14912 17380 14916 17436
rect 14852 17376 14916 17380
rect 14932 17436 14996 17440
rect 14932 17380 14936 17436
rect 14936 17380 14992 17436
rect 14992 17380 14996 17436
rect 14932 17376 14996 17380
rect 15012 17436 15076 17440
rect 15012 17380 15016 17436
rect 15016 17380 15072 17436
rect 15072 17380 15076 17436
rect 15012 17376 15076 17380
rect 15092 17436 15156 17440
rect 15092 17380 15096 17436
rect 15096 17380 15152 17436
rect 15152 17380 15156 17436
rect 15092 17376 15156 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 17932 17436 17996 17440
rect 17932 17380 17936 17436
rect 17936 17380 17992 17436
rect 17992 17380 17996 17436
rect 17932 17376 17996 17380
rect 18012 17436 18076 17440
rect 18012 17380 18016 17436
rect 18016 17380 18072 17436
rect 18072 17380 18076 17436
rect 18012 17376 18076 17380
rect 18092 17436 18156 17440
rect 18092 17380 18096 17436
rect 18096 17380 18152 17436
rect 18152 17380 18156 17436
rect 18092 17376 18156 17380
rect 20852 17436 20916 17440
rect 20852 17380 20856 17436
rect 20856 17380 20912 17436
rect 20912 17380 20916 17436
rect 20852 17376 20916 17380
rect 20932 17436 20996 17440
rect 20932 17380 20936 17436
rect 20936 17380 20992 17436
rect 20992 17380 20996 17436
rect 20932 17376 20996 17380
rect 21012 17436 21076 17440
rect 21012 17380 21016 17436
rect 21016 17380 21072 17436
rect 21072 17380 21076 17436
rect 21012 17376 21076 17380
rect 21092 17436 21156 17440
rect 21092 17380 21096 17436
rect 21096 17380 21152 17436
rect 21152 17380 21156 17436
rect 21092 17376 21156 17380
rect 23852 17436 23916 17440
rect 23852 17380 23856 17436
rect 23856 17380 23912 17436
rect 23912 17380 23916 17436
rect 23852 17376 23916 17380
rect 23932 17436 23996 17440
rect 23932 17380 23936 17436
rect 23936 17380 23992 17436
rect 23992 17380 23996 17436
rect 23932 17376 23996 17380
rect 24012 17436 24076 17440
rect 24012 17380 24016 17436
rect 24016 17380 24072 17436
rect 24072 17380 24076 17436
rect 24012 17376 24076 17380
rect 24092 17436 24156 17440
rect 24092 17380 24096 17436
rect 24096 17380 24152 17436
rect 24152 17380 24156 17436
rect 24092 17376 24156 17380
rect 1352 16892 1416 16896
rect 1352 16836 1356 16892
rect 1356 16836 1412 16892
rect 1412 16836 1416 16892
rect 1352 16832 1416 16836
rect 1432 16892 1496 16896
rect 1432 16836 1436 16892
rect 1436 16836 1492 16892
rect 1492 16836 1496 16892
rect 1432 16832 1496 16836
rect 1512 16892 1576 16896
rect 1512 16836 1516 16892
rect 1516 16836 1572 16892
rect 1572 16836 1576 16892
rect 1512 16832 1576 16836
rect 1592 16892 1656 16896
rect 1592 16836 1596 16892
rect 1596 16836 1652 16892
rect 1652 16836 1656 16892
rect 1592 16832 1656 16836
rect 4352 16892 4416 16896
rect 4352 16836 4356 16892
rect 4356 16836 4412 16892
rect 4412 16836 4416 16892
rect 4352 16832 4416 16836
rect 4432 16892 4496 16896
rect 4432 16836 4436 16892
rect 4436 16836 4492 16892
rect 4492 16836 4496 16892
rect 4432 16832 4496 16836
rect 4512 16892 4576 16896
rect 4512 16836 4516 16892
rect 4516 16836 4572 16892
rect 4572 16836 4576 16892
rect 4512 16832 4576 16836
rect 4592 16892 4656 16896
rect 4592 16836 4596 16892
rect 4596 16836 4652 16892
rect 4652 16836 4656 16892
rect 4592 16832 4656 16836
rect 7352 16892 7416 16896
rect 7352 16836 7356 16892
rect 7356 16836 7412 16892
rect 7412 16836 7416 16892
rect 7352 16832 7416 16836
rect 7432 16892 7496 16896
rect 7432 16836 7436 16892
rect 7436 16836 7492 16892
rect 7492 16836 7496 16892
rect 7432 16832 7496 16836
rect 7512 16892 7576 16896
rect 7512 16836 7516 16892
rect 7516 16836 7572 16892
rect 7572 16836 7576 16892
rect 7512 16832 7576 16836
rect 7592 16892 7656 16896
rect 7592 16836 7596 16892
rect 7596 16836 7652 16892
rect 7652 16836 7656 16892
rect 7592 16832 7656 16836
rect 10352 16892 10416 16896
rect 10352 16836 10356 16892
rect 10356 16836 10412 16892
rect 10412 16836 10416 16892
rect 10352 16832 10416 16836
rect 10432 16892 10496 16896
rect 10432 16836 10436 16892
rect 10436 16836 10492 16892
rect 10492 16836 10496 16892
rect 10432 16832 10496 16836
rect 10512 16892 10576 16896
rect 10512 16836 10516 16892
rect 10516 16836 10572 16892
rect 10572 16836 10576 16892
rect 10512 16832 10576 16836
rect 10592 16892 10656 16896
rect 10592 16836 10596 16892
rect 10596 16836 10652 16892
rect 10652 16836 10656 16892
rect 10592 16832 10656 16836
rect 13352 16892 13416 16896
rect 13352 16836 13356 16892
rect 13356 16836 13412 16892
rect 13412 16836 13416 16892
rect 13352 16832 13416 16836
rect 13432 16892 13496 16896
rect 13432 16836 13436 16892
rect 13436 16836 13492 16892
rect 13492 16836 13496 16892
rect 13432 16832 13496 16836
rect 13512 16892 13576 16896
rect 13512 16836 13516 16892
rect 13516 16836 13572 16892
rect 13572 16836 13576 16892
rect 13512 16832 13576 16836
rect 13592 16892 13656 16896
rect 13592 16836 13596 16892
rect 13596 16836 13652 16892
rect 13652 16836 13656 16892
rect 13592 16832 13656 16836
rect 16352 16892 16416 16896
rect 16352 16836 16356 16892
rect 16356 16836 16412 16892
rect 16412 16836 16416 16892
rect 16352 16832 16416 16836
rect 16432 16892 16496 16896
rect 16432 16836 16436 16892
rect 16436 16836 16492 16892
rect 16492 16836 16496 16892
rect 16432 16832 16496 16836
rect 16512 16892 16576 16896
rect 16512 16836 16516 16892
rect 16516 16836 16572 16892
rect 16572 16836 16576 16892
rect 16512 16832 16576 16836
rect 16592 16892 16656 16896
rect 16592 16836 16596 16892
rect 16596 16836 16652 16892
rect 16652 16836 16656 16892
rect 16592 16832 16656 16836
rect 19352 16892 19416 16896
rect 19352 16836 19356 16892
rect 19356 16836 19412 16892
rect 19412 16836 19416 16892
rect 19352 16832 19416 16836
rect 19432 16892 19496 16896
rect 19432 16836 19436 16892
rect 19436 16836 19492 16892
rect 19492 16836 19496 16892
rect 19432 16832 19496 16836
rect 19512 16892 19576 16896
rect 19512 16836 19516 16892
rect 19516 16836 19572 16892
rect 19572 16836 19576 16892
rect 19512 16832 19576 16836
rect 19592 16892 19656 16896
rect 19592 16836 19596 16892
rect 19596 16836 19652 16892
rect 19652 16836 19656 16892
rect 19592 16832 19656 16836
rect 22352 16892 22416 16896
rect 22352 16836 22356 16892
rect 22356 16836 22412 16892
rect 22412 16836 22416 16892
rect 22352 16832 22416 16836
rect 22432 16892 22496 16896
rect 22432 16836 22436 16892
rect 22436 16836 22492 16892
rect 22492 16836 22496 16892
rect 22432 16832 22496 16836
rect 22512 16892 22576 16896
rect 22512 16836 22516 16892
rect 22516 16836 22572 16892
rect 22572 16836 22576 16892
rect 22512 16832 22576 16836
rect 22592 16892 22656 16896
rect 22592 16836 22596 16892
rect 22596 16836 22652 16892
rect 22652 16836 22656 16892
rect 22592 16832 22656 16836
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 2932 16348 2996 16352
rect 2932 16292 2936 16348
rect 2936 16292 2992 16348
rect 2992 16292 2996 16348
rect 2932 16288 2996 16292
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 5852 16348 5916 16352
rect 5852 16292 5856 16348
rect 5856 16292 5912 16348
rect 5912 16292 5916 16348
rect 5852 16288 5916 16292
rect 5932 16348 5996 16352
rect 5932 16292 5936 16348
rect 5936 16292 5992 16348
rect 5992 16292 5996 16348
rect 5932 16288 5996 16292
rect 6012 16348 6076 16352
rect 6012 16292 6016 16348
rect 6016 16292 6072 16348
rect 6072 16292 6076 16348
rect 6012 16288 6076 16292
rect 6092 16348 6156 16352
rect 6092 16292 6096 16348
rect 6096 16292 6152 16348
rect 6152 16292 6156 16348
rect 6092 16288 6156 16292
rect 8852 16348 8916 16352
rect 8852 16292 8856 16348
rect 8856 16292 8912 16348
rect 8912 16292 8916 16348
rect 8852 16288 8916 16292
rect 8932 16348 8996 16352
rect 8932 16292 8936 16348
rect 8936 16292 8992 16348
rect 8992 16292 8996 16348
rect 8932 16288 8996 16292
rect 9012 16348 9076 16352
rect 9012 16292 9016 16348
rect 9016 16292 9072 16348
rect 9072 16292 9076 16348
rect 9012 16288 9076 16292
rect 9092 16348 9156 16352
rect 9092 16292 9096 16348
rect 9096 16292 9152 16348
rect 9152 16292 9156 16348
rect 9092 16288 9156 16292
rect 11852 16348 11916 16352
rect 11852 16292 11856 16348
rect 11856 16292 11912 16348
rect 11912 16292 11916 16348
rect 11852 16288 11916 16292
rect 11932 16348 11996 16352
rect 11932 16292 11936 16348
rect 11936 16292 11992 16348
rect 11992 16292 11996 16348
rect 11932 16288 11996 16292
rect 12012 16348 12076 16352
rect 12012 16292 12016 16348
rect 12016 16292 12072 16348
rect 12072 16292 12076 16348
rect 12012 16288 12076 16292
rect 12092 16348 12156 16352
rect 12092 16292 12096 16348
rect 12096 16292 12152 16348
rect 12152 16292 12156 16348
rect 12092 16288 12156 16292
rect 14852 16348 14916 16352
rect 14852 16292 14856 16348
rect 14856 16292 14912 16348
rect 14912 16292 14916 16348
rect 14852 16288 14916 16292
rect 14932 16348 14996 16352
rect 14932 16292 14936 16348
rect 14936 16292 14992 16348
rect 14992 16292 14996 16348
rect 14932 16288 14996 16292
rect 15012 16348 15076 16352
rect 15012 16292 15016 16348
rect 15016 16292 15072 16348
rect 15072 16292 15076 16348
rect 15012 16288 15076 16292
rect 15092 16348 15156 16352
rect 15092 16292 15096 16348
rect 15096 16292 15152 16348
rect 15152 16292 15156 16348
rect 15092 16288 15156 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 17932 16348 17996 16352
rect 17932 16292 17936 16348
rect 17936 16292 17992 16348
rect 17992 16292 17996 16348
rect 17932 16288 17996 16292
rect 18012 16348 18076 16352
rect 18012 16292 18016 16348
rect 18016 16292 18072 16348
rect 18072 16292 18076 16348
rect 18012 16288 18076 16292
rect 18092 16348 18156 16352
rect 18092 16292 18096 16348
rect 18096 16292 18152 16348
rect 18152 16292 18156 16348
rect 18092 16288 18156 16292
rect 20852 16348 20916 16352
rect 20852 16292 20856 16348
rect 20856 16292 20912 16348
rect 20912 16292 20916 16348
rect 20852 16288 20916 16292
rect 20932 16348 20996 16352
rect 20932 16292 20936 16348
rect 20936 16292 20992 16348
rect 20992 16292 20996 16348
rect 20932 16288 20996 16292
rect 21012 16348 21076 16352
rect 21012 16292 21016 16348
rect 21016 16292 21072 16348
rect 21072 16292 21076 16348
rect 21012 16288 21076 16292
rect 21092 16348 21156 16352
rect 21092 16292 21096 16348
rect 21096 16292 21152 16348
rect 21152 16292 21156 16348
rect 21092 16288 21156 16292
rect 23852 16348 23916 16352
rect 23852 16292 23856 16348
rect 23856 16292 23912 16348
rect 23912 16292 23916 16348
rect 23852 16288 23916 16292
rect 23932 16348 23996 16352
rect 23932 16292 23936 16348
rect 23936 16292 23992 16348
rect 23992 16292 23996 16348
rect 23932 16288 23996 16292
rect 24012 16348 24076 16352
rect 24012 16292 24016 16348
rect 24016 16292 24072 16348
rect 24072 16292 24076 16348
rect 24012 16288 24076 16292
rect 24092 16348 24156 16352
rect 24092 16292 24096 16348
rect 24096 16292 24152 16348
rect 24152 16292 24156 16348
rect 24092 16288 24156 16292
rect 1352 15804 1416 15808
rect 1352 15748 1356 15804
rect 1356 15748 1412 15804
rect 1412 15748 1416 15804
rect 1352 15744 1416 15748
rect 1432 15804 1496 15808
rect 1432 15748 1436 15804
rect 1436 15748 1492 15804
rect 1492 15748 1496 15804
rect 1432 15744 1496 15748
rect 1512 15804 1576 15808
rect 1512 15748 1516 15804
rect 1516 15748 1572 15804
rect 1572 15748 1576 15804
rect 1512 15744 1576 15748
rect 1592 15804 1656 15808
rect 1592 15748 1596 15804
rect 1596 15748 1652 15804
rect 1652 15748 1656 15804
rect 1592 15744 1656 15748
rect 4352 15804 4416 15808
rect 4352 15748 4356 15804
rect 4356 15748 4412 15804
rect 4412 15748 4416 15804
rect 4352 15744 4416 15748
rect 4432 15804 4496 15808
rect 4432 15748 4436 15804
rect 4436 15748 4492 15804
rect 4492 15748 4496 15804
rect 4432 15744 4496 15748
rect 4512 15804 4576 15808
rect 4512 15748 4516 15804
rect 4516 15748 4572 15804
rect 4572 15748 4576 15804
rect 4512 15744 4576 15748
rect 4592 15804 4656 15808
rect 4592 15748 4596 15804
rect 4596 15748 4652 15804
rect 4652 15748 4656 15804
rect 4592 15744 4656 15748
rect 7352 15804 7416 15808
rect 7352 15748 7356 15804
rect 7356 15748 7412 15804
rect 7412 15748 7416 15804
rect 7352 15744 7416 15748
rect 7432 15804 7496 15808
rect 7432 15748 7436 15804
rect 7436 15748 7492 15804
rect 7492 15748 7496 15804
rect 7432 15744 7496 15748
rect 7512 15804 7576 15808
rect 7512 15748 7516 15804
rect 7516 15748 7572 15804
rect 7572 15748 7576 15804
rect 7512 15744 7576 15748
rect 7592 15804 7656 15808
rect 7592 15748 7596 15804
rect 7596 15748 7652 15804
rect 7652 15748 7656 15804
rect 7592 15744 7656 15748
rect 10352 15804 10416 15808
rect 10352 15748 10356 15804
rect 10356 15748 10412 15804
rect 10412 15748 10416 15804
rect 10352 15744 10416 15748
rect 10432 15804 10496 15808
rect 10432 15748 10436 15804
rect 10436 15748 10492 15804
rect 10492 15748 10496 15804
rect 10432 15744 10496 15748
rect 10512 15804 10576 15808
rect 10512 15748 10516 15804
rect 10516 15748 10572 15804
rect 10572 15748 10576 15804
rect 10512 15744 10576 15748
rect 10592 15804 10656 15808
rect 10592 15748 10596 15804
rect 10596 15748 10652 15804
rect 10652 15748 10656 15804
rect 10592 15744 10656 15748
rect 13352 15804 13416 15808
rect 13352 15748 13356 15804
rect 13356 15748 13412 15804
rect 13412 15748 13416 15804
rect 13352 15744 13416 15748
rect 13432 15804 13496 15808
rect 13432 15748 13436 15804
rect 13436 15748 13492 15804
rect 13492 15748 13496 15804
rect 13432 15744 13496 15748
rect 13512 15804 13576 15808
rect 13512 15748 13516 15804
rect 13516 15748 13572 15804
rect 13572 15748 13576 15804
rect 13512 15744 13576 15748
rect 13592 15804 13656 15808
rect 13592 15748 13596 15804
rect 13596 15748 13652 15804
rect 13652 15748 13656 15804
rect 13592 15744 13656 15748
rect 16352 15804 16416 15808
rect 16352 15748 16356 15804
rect 16356 15748 16412 15804
rect 16412 15748 16416 15804
rect 16352 15744 16416 15748
rect 16432 15804 16496 15808
rect 16432 15748 16436 15804
rect 16436 15748 16492 15804
rect 16492 15748 16496 15804
rect 16432 15744 16496 15748
rect 16512 15804 16576 15808
rect 16512 15748 16516 15804
rect 16516 15748 16572 15804
rect 16572 15748 16576 15804
rect 16512 15744 16576 15748
rect 16592 15804 16656 15808
rect 16592 15748 16596 15804
rect 16596 15748 16652 15804
rect 16652 15748 16656 15804
rect 16592 15744 16656 15748
rect 19352 15804 19416 15808
rect 19352 15748 19356 15804
rect 19356 15748 19412 15804
rect 19412 15748 19416 15804
rect 19352 15744 19416 15748
rect 19432 15804 19496 15808
rect 19432 15748 19436 15804
rect 19436 15748 19492 15804
rect 19492 15748 19496 15804
rect 19432 15744 19496 15748
rect 19512 15804 19576 15808
rect 19512 15748 19516 15804
rect 19516 15748 19572 15804
rect 19572 15748 19576 15804
rect 19512 15744 19576 15748
rect 19592 15804 19656 15808
rect 19592 15748 19596 15804
rect 19596 15748 19652 15804
rect 19652 15748 19656 15804
rect 19592 15744 19656 15748
rect 22352 15804 22416 15808
rect 22352 15748 22356 15804
rect 22356 15748 22412 15804
rect 22412 15748 22416 15804
rect 22352 15744 22416 15748
rect 22432 15804 22496 15808
rect 22432 15748 22436 15804
rect 22436 15748 22492 15804
rect 22492 15748 22496 15804
rect 22432 15744 22496 15748
rect 22512 15804 22576 15808
rect 22512 15748 22516 15804
rect 22516 15748 22572 15804
rect 22572 15748 22576 15804
rect 22512 15744 22576 15748
rect 22592 15804 22656 15808
rect 22592 15748 22596 15804
rect 22596 15748 22652 15804
rect 22652 15748 22656 15804
rect 22592 15744 22656 15748
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 2932 15260 2996 15264
rect 2932 15204 2936 15260
rect 2936 15204 2992 15260
rect 2992 15204 2996 15260
rect 2932 15200 2996 15204
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 5852 15260 5916 15264
rect 5852 15204 5856 15260
rect 5856 15204 5912 15260
rect 5912 15204 5916 15260
rect 5852 15200 5916 15204
rect 5932 15260 5996 15264
rect 5932 15204 5936 15260
rect 5936 15204 5992 15260
rect 5992 15204 5996 15260
rect 5932 15200 5996 15204
rect 6012 15260 6076 15264
rect 6012 15204 6016 15260
rect 6016 15204 6072 15260
rect 6072 15204 6076 15260
rect 6012 15200 6076 15204
rect 6092 15260 6156 15264
rect 6092 15204 6096 15260
rect 6096 15204 6152 15260
rect 6152 15204 6156 15260
rect 6092 15200 6156 15204
rect 8852 15260 8916 15264
rect 8852 15204 8856 15260
rect 8856 15204 8912 15260
rect 8912 15204 8916 15260
rect 8852 15200 8916 15204
rect 8932 15260 8996 15264
rect 8932 15204 8936 15260
rect 8936 15204 8992 15260
rect 8992 15204 8996 15260
rect 8932 15200 8996 15204
rect 9012 15260 9076 15264
rect 9012 15204 9016 15260
rect 9016 15204 9072 15260
rect 9072 15204 9076 15260
rect 9012 15200 9076 15204
rect 9092 15260 9156 15264
rect 9092 15204 9096 15260
rect 9096 15204 9152 15260
rect 9152 15204 9156 15260
rect 9092 15200 9156 15204
rect 11852 15260 11916 15264
rect 11852 15204 11856 15260
rect 11856 15204 11912 15260
rect 11912 15204 11916 15260
rect 11852 15200 11916 15204
rect 11932 15260 11996 15264
rect 11932 15204 11936 15260
rect 11936 15204 11992 15260
rect 11992 15204 11996 15260
rect 11932 15200 11996 15204
rect 12012 15260 12076 15264
rect 12012 15204 12016 15260
rect 12016 15204 12072 15260
rect 12072 15204 12076 15260
rect 12012 15200 12076 15204
rect 12092 15260 12156 15264
rect 12092 15204 12096 15260
rect 12096 15204 12152 15260
rect 12152 15204 12156 15260
rect 12092 15200 12156 15204
rect 14852 15260 14916 15264
rect 14852 15204 14856 15260
rect 14856 15204 14912 15260
rect 14912 15204 14916 15260
rect 14852 15200 14916 15204
rect 14932 15260 14996 15264
rect 14932 15204 14936 15260
rect 14936 15204 14992 15260
rect 14992 15204 14996 15260
rect 14932 15200 14996 15204
rect 15012 15260 15076 15264
rect 15012 15204 15016 15260
rect 15016 15204 15072 15260
rect 15072 15204 15076 15260
rect 15012 15200 15076 15204
rect 15092 15260 15156 15264
rect 15092 15204 15096 15260
rect 15096 15204 15152 15260
rect 15152 15204 15156 15260
rect 15092 15200 15156 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 17932 15260 17996 15264
rect 17932 15204 17936 15260
rect 17936 15204 17992 15260
rect 17992 15204 17996 15260
rect 17932 15200 17996 15204
rect 18012 15260 18076 15264
rect 18012 15204 18016 15260
rect 18016 15204 18072 15260
rect 18072 15204 18076 15260
rect 18012 15200 18076 15204
rect 18092 15260 18156 15264
rect 18092 15204 18096 15260
rect 18096 15204 18152 15260
rect 18152 15204 18156 15260
rect 18092 15200 18156 15204
rect 20852 15260 20916 15264
rect 20852 15204 20856 15260
rect 20856 15204 20912 15260
rect 20912 15204 20916 15260
rect 20852 15200 20916 15204
rect 20932 15260 20996 15264
rect 20932 15204 20936 15260
rect 20936 15204 20992 15260
rect 20992 15204 20996 15260
rect 20932 15200 20996 15204
rect 21012 15260 21076 15264
rect 21012 15204 21016 15260
rect 21016 15204 21072 15260
rect 21072 15204 21076 15260
rect 21012 15200 21076 15204
rect 21092 15260 21156 15264
rect 21092 15204 21096 15260
rect 21096 15204 21152 15260
rect 21152 15204 21156 15260
rect 21092 15200 21156 15204
rect 23852 15260 23916 15264
rect 23852 15204 23856 15260
rect 23856 15204 23912 15260
rect 23912 15204 23916 15260
rect 23852 15200 23916 15204
rect 23932 15260 23996 15264
rect 23932 15204 23936 15260
rect 23936 15204 23992 15260
rect 23992 15204 23996 15260
rect 23932 15200 23996 15204
rect 24012 15260 24076 15264
rect 24012 15204 24016 15260
rect 24016 15204 24072 15260
rect 24072 15204 24076 15260
rect 24012 15200 24076 15204
rect 24092 15260 24156 15264
rect 24092 15204 24096 15260
rect 24096 15204 24152 15260
rect 24152 15204 24156 15260
rect 24092 15200 24156 15204
rect 1352 14716 1416 14720
rect 1352 14660 1356 14716
rect 1356 14660 1412 14716
rect 1412 14660 1416 14716
rect 1352 14656 1416 14660
rect 1432 14716 1496 14720
rect 1432 14660 1436 14716
rect 1436 14660 1492 14716
rect 1492 14660 1496 14716
rect 1432 14656 1496 14660
rect 1512 14716 1576 14720
rect 1512 14660 1516 14716
rect 1516 14660 1572 14716
rect 1572 14660 1576 14716
rect 1512 14656 1576 14660
rect 1592 14716 1656 14720
rect 1592 14660 1596 14716
rect 1596 14660 1652 14716
rect 1652 14660 1656 14716
rect 1592 14656 1656 14660
rect 4352 14716 4416 14720
rect 4352 14660 4356 14716
rect 4356 14660 4412 14716
rect 4412 14660 4416 14716
rect 4352 14656 4416 14660
rect 4432 14716 4496 14720
rect 4432 14660 4436 14716
rect 4436 14660 4492 14716
rect 4492 14660 4496 14716
rect 4432 14656 4496 14660
rect 4512 14716 4576 14720
rect 4512 14660 4516 14716
rect 4516 14660 4572 14716
rect 4572 14660 4576 14716
rect 4512 14656 4576 14660
rect 4592 14716 4656 14720
rect 4592 14660 4596 14716
rect 4596 14660 4652 14716
rect 4652 14660 4656 14716
rect 4592 14656 4656 14660
rect 7352 14716 7416 14720
rect 7352 14660 7356 14716
rect 7356 14660 7412 14716
rect 7412 14660 7416 14716
rect 7352 14656 7416 14660
rect 7432 14716 7496 14720
rect 7432 14660 7436 14716
rect 7436 14660 7492 14716
rect 7492 14660 7496 14716
rect 7432 14656 7496 14660
rect 7512 14716 7576 14720
rect 7512 14660 7516 14716
rect 7516 14660 7572 14716
rect 7572 14660 7576 14716
rect 7512 14656 7576 14660
rect 7592 14716 7656 14720
rect 7592 14660 7596 14716
rect 7596 14660 7652 14716
rect 7652 14660 7656 14716
rect 7592 14656 7656 14660
rect 10352 14716 10416 14720
rect 10352 14660 10356 14716
rect 10356 14660 10412 14716
rect 10412 14660 10416 14716
rect 10352 14656 10416 14660
rect 10432 14716 10496 14720
rect 10432 14660 10436 14716
rect 10436 14660 10492 14716
rect 10492 14660 10496 14716
rect 10432 14656 10496 14660
rect 10512 14716 10576 14720
rect 10512 14660 10516 14716
rect 10516 14660 10572 14716
rect 10572 14660 10576 14716
rect 10512 14656 10576 14660
rect 10592 14716 10656 14720
rect 10592 14660 10596 14716
rect 10596 14660 10652 14716
rect 10652 14660 10656 14716
rect 10592 14656 10656 14660
rect 13352 14716 13416 14720
rect 13352 14660 13356 14716
rect 13356 14660 13412 14716
rect 13412 14660 13416 14716
rect 13352 14656 13416 14660
rect 13432 14716 13496 14720
rect 13432 14660 13436 14716
rect 13436 14660 13492 14716
rect 13492 14660 13496 14716
rect 13432 14656 13496 14660
rect 13512 14716 13576 14720
rect 13512 14660 13516 14716
rect 13516 14660 13572 14716
rect 13572 14660 13576 14716
rect 13512 14656 13576 14660
rect 13592 14716 13656 14720
rect 13592 14660 13596 14716
rect 13596 14660 13652 14716
rect 13652 14660 13656 14716
rect 13592 14656 13656 14660
rect 16352 14716 16416 14720
rect 16352 14660 16356 14716
rect 16356 14660 16412 14716
rect 16412 14660 16416 14716
rect 16352 14656 16416 14660
rect 16432 14716 16496 14720
rect 16432 14660 16436 14716
rect 16436 14660 16492 14716
rect 16492 14660 16496 14716
rect 16432 14656 16496 14660
rect 16512 14716 16576 14720
rect 16512 14660 16516 14716
rect 16516 14660 16572 14716
rect 16572 14660 16576 14716
rect 16512 14656 16576 14660
rect 16592 14716 16656 14720
rect 16592 14660 16596 14716
rect 16596 14660 16652 14716
rect 16652 14660 16656 14716
rect 16592 14656 16656 14660
rect 19352 14716 19416 14720
rect 19352 14660 19356 14716
rect 19356 14660 19412 14716
rect 19412 14660 19416 14716
rect 19352 14656 19416 14660
rect 19432 14716 19496 14720
rect 19432 14660 19436 14716
rect 19436 14660 19492 14716
rect 19492 14660 19496 14716
rect 19432 14656 19496 14660
rect 19512 14716 19576 14720
rect 19512 14660 19516 14716
rect 19516 14660 19572 14716
rect 19572 14660 19576 14716
rect 19512 14656 19576 14660
rect 19592 14716 19656 14720
rect 19592 14660 19596 14716
rect 19596 14660 19652 14716
rect 19652 14660 19656 14716
rect 19592 14656 19656 14660
rect 22352 14716 22416 14720
rect 22352 14660 22356 14716
rect 22356 14660 22412 14716
rect 22412 14660 22416 14716
rect 22352 14656 22416 14660
rect 22432 14716 22496 14720
rect 22432 14660 22436 14716
rect 22436 14660 22492 14716
rect 22492 14660 22496 14716
rect 22432 14656 22496 14660
rect 22512 14716 22576 14720
rect 22512 14660 22516 14716
rect 22516 14660 22572 14716
rect 22572 14660 22576 14716
rect 22512 14656 22576 14660
rect 22592 14716 22656 14720
rect 22592 14660 22596 14716
rect 22596 14660 22652 14716
rect 22652 14660 22656 14716
rect 22592 14656 22656 14660
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 2932 14172 2996 14176
rect 2932 14116 2936 14172
rect 2936 14116 2992 14172
rect 2992 14116 2996 14172
rect 2932 14112 2996 14116
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 5852 14172 5916 14176
rect 5852 14116 5856 14172
rect 5856 14116 5912 14172
rect 5912 14116 5916 14172
rect 5852 14112 5916 14116
rect 5932 14172 5996 14176
rect 5932 14116 5936 14172
rect 5936 14116 5992 14172
rect 5992 14116 5996 14172
rect 5932 14112 5996 14116
rect 6012 14172 6076 14176
rect 6012 14116 6016 14172
rect 6016 14116 6072 14172
rect 6072 14116 6076 14172
rect 6012 14112 6076 14116
rect 6092 14172 6156 14176
rect 6092 14116 6096 14172
rect 6096 14116 6152 14172
rect 6152 14116 6156 14172
rect 6092 14112 6156 14116
rect 8852 14172 8916 14176
rect 8852 14116 8856 14172
rect 8856 14116 8912 14172
rect 8912 14116 8916 14172
rect 8852 14112 8916 14116
rect 8932 14172 8996 14176
rect 8932 14116 8936 14172
rect 8936 14116 8992 14172
rect 8992 14116 8996 14172
rect 8932 14112 8996 14116
rect 9012 14172 9076 14176
rect 9012 14116 9016 14172
rect 9016 14116 9072 14172
rect 9072 14116 9076 14172
rect 9012 14112 9076 14116
rect 9092 14172 9156 14176
rect 9092 14116 9096 14172
rect 9096 14116 9152 14172
rect 9152 14116 9156 14172
rect 9092 14112 9156 14116
rect 11852 14172 11916 14176
rect 11852 14116 11856 14172
rect 11856 14116 11912 14172
rect 11912 14116 11916 14172
rect 11852 14112 11916 14116
rect 11932 14172 11996 14176
rect 11932 14116 11936 14172
rect 11936 14116 11992 14172
rect 11992 14116 11996 14172
rect 11932 14112 11996 14116
rect 12012 14172 12076 14176
rect 12012 14116 12016 14172
rect 12016 14116 12072 14172
rect 12072 14116 12076 14172
rect 12012 14112 12076 14116
rect 12092 14172 12156 14176
rect 12092 14116 12096 14172
rect 12096 14116 12152 14172
rect 12152 14116 12156 14172
rect 12092 14112 12156 14116
rect 14852 14172 14916 14176
rect 14852 14116 14856 14172
rect 14856 14116 14912 14172
rect 14912 14116 14916 14172
rect 14852 14112 14916 14116
rect 14932 14172 14996 14176
rect 14932 14116 14936 14172
rect 14936 14116 14992 14172
rect 14992 14116 14996 14172
rect 14932 14112 14996 14116
rect 15012 14172 15076 14176
rect 15012 14116 15016 14172
rect 15016 14116 15072 14172
rect 15072 14116 15076 14172
rect 15012 14112 15076 14116
rect 15092 14172 15156 14176
rect 15092 14116 15096 14172
rect 15096 14116 15152 14172
rect 15152 14116 15156 14172
rect 15092 14112 15156 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 17932 14172 17996 14176
rect 17932 14116 17936 14172
rect 17936 14116 17992 14172
rect 17992 14116 17996 14172
rect 17932 14112 17996 14116
rect 18012 14172 18076 14176
rect 18012 14116 18016 14172
rect 18016 14116 18072 14172
rect 18072 14116 18076 14172
rect 18012 14112 18076 14116
rect 18092 14172 18156 14176
rect 18092 14116 18096 14172
rect 18096 14116 18152 14172
rect 18152 14116 18156 14172
rect 18092 14112 18156 14116
rect 20852 14172 20916 14176
rect 20852 14116 20856 14172
rect 20856 14116 20912 14172
rect 20912 14116 20916 14172
rect 20852 14112 20916 14116
rect 20932 14172 20996 14176
rect 20932 14116 20936 14172
rect 20936 14116 20992 14172
rect 20992 14116 20996 14172
rect 20932 14112 20996 14116
rect 21012 14172 21076 14176
rect 21012 14116 21016 14172
rect 21016 14116 21072 14172
rect 21072 14116 21076 14172
rect 21012 14112 21076 14116
rect 21092 14172 21156 14176
rect 21092 14116 21096 14172
rect 21096 14116 21152 14172
rect 21152 14116 21156 14172
rect 21092 14112 21156 14116
rect 23852 14172 23916 14176
rect 23852 14116 23856 14172
rect 23856 14116 23912 14172
rect 23912 14116 23916 14172
rect 23852 14112 23916 14116
rect 23932 14172 23996 14176
rect 23932 14116 23936 14172
rect 23936 14116 23992 14172
rect 23992 14116 23996 14172
rect 23932 14112 23996 14116
rect 24012 14172 24076 14176
rect 24012 14116 24016 14172
rect 24016 14116 24072 14172
rect 24072 14116 24076 14172
rect 24012 14112 24076 14116
rect 24092 14172 24156 14176
rect 24092 14116 24096 14172
rect 24096 14116 24152 14172
rect 24152 14116 24156 14172
rect 24092 14112 24156 14116
rect 3372 13908 3436 13972
rect 13124 13908 13188 13972
rect 22140 13696 22204 13700
rect 22140 13640 22154 13696
rect 22154 13640 22204 13696
rect 22140 13636 22204 13640
rect 1352 13628 1416 13632
rect 1352 13572 1356 13628
rect 1356 13572 1412 13628
rect 1412 13572 1416 13628
rect 1352 13568 1416 13572
rect 1432 13628 1496 13632
rect 1432 13572 1436 13628
rect 1436 13572 1492 13628
rect 1492 13572 1496 13628
rect 1432 13568 1496 13572
rect 1512 13628 1576 13632
rect 1512 13572 1516 13628
rect 1516 13572 1572 13628
rect 1572 13572 1576 13628
rect 1512 13568 1576 13572
rect 1592 13628 1656 13632
rect 1592 13572 1596 13628
rect 1596 13572 1652 13628
rect 1652 13572 1656 13628
rect 1592 13568 1656 13572
rect 4352 13628 4416 13632
rect 4352 13572 4356 13628
rect 4356 13572 4412 13628
rect 4412 13572 4416 13628
rect 4352 13568 4416 13572
rect 4432 13628 4496 13632
rect 4432 13572 4436 13628
rect 4436 13572 4492 13628
rect 4492 13572 4496 13628
rect 4432 13568 4496 13572
rect 4512 13628 4576 13632
rect 4512 13572 4516 13628
rect 4516 13572 4572 13628
rect 4572 13572 4576 13628
rect 4512 13568 4576 13572
rect 4592 13628 4656 13632
rect 4592 13572 4596 13628
rect 4596 13572 4652 13628
rect 4652 13572 4656 13628
rect 4592 13568 4656 13572
rect 7352 13628 7416 13632
rect 7352 13572 7356 13628
rect 7356 13572 7412 13628
rect 7412 13572 7416 13628
rect 7352 13568 7416 13572
rect 7432 13628 7496 13632
rect 7432 13572 7436 13628
rect 7436 13572 7492 13628
rect 7492 13572 7496 13628
rect 7432 13568 7496 13572
rect 7512 13628 7576 13632
rect 7512 13572 7516 13628
rect 7516 13572 7572 13628
rect 7572 13572 7576 13628
rect 7512 13568 7576 13572
rect 7592 13628 7656 13632
rect 7592 13572 7596 13628
rect 7596 13572 7652 13628
rect 7652 13572 7656 13628
rect 7592 13568 7656 13572
rect 10352 13628 10416 13632
rect 10352 13572 10356 13628
rect 10356 13572 10412 13628
rect 10412 13572 10416 13628
rect 10352 13568 10416 13572
rect 10432 13628 10496 13632
rect 10432 13572 10436 13628
rect 10436 13572 10492 13628
rect 10492 13572 10496 13628
rect 10432 13568 10496 13572
rect 10512 13628 10576 13632
rect 10512 13572 10516 13628
rect 10516 13572 10572 13628
rect 10572 13572 10576 13628
rect 10512 13568 10576 13572
rect 10592 13628 10656 13632
rect 10592 13572 10596 13628
rect 10596 13572 10652 13628
rect 10652 13572 10656 13628
rect 10592 13568 10656 13572
rect 13352 13628 13416 13632
rect 13352 13572 13356 13628
rect 13356 13572 13412 13628
rect 13412 13572 13416 13628
rect 13352 13568 13416 13572
rect 13432 13628 13496 13632
rect 13432 13572 13436 13628
rect 13436 13572 13492 13628
rect 13492 13572 13496 13628
rect 13432 13568 13496 13572
rect 13512 13628 13576 13632
rect 13512 13572 13516 13628
rect 13516 13572 13572 13628
rect 13572 13572 13576 13628
rect 13512 13568 13576 13572
rect 13592 13628 13656 13632
rect 13592 13572 13596 13628
rect 13596 13572 13652 13628
rect 13652 13572 13656 13628
rect 13592 13568 13656 13572
rect 16352 13628 16416 13632
rect 16352 13572 16356 13628
rect 16356 13572 16412 13628
rect 16412 13572 16416 13628
rect 16352 13568 16416 13572
rect 16432 13628 16496 13632
rect 16432 13572 16436 13628
rect 16436 13572 16492 13628
rect 16492 13572 16496 13628
rect 16432 13568 16496 13572
rect 16512 13628 16576 13632
rect 16512 13572 16516 13628
rect 16516 13572 16572 13628
rect 16572 13572 16576 13628
rect 16512 13568 16576 13572
rect 16592 13628 16656 13632
rect 16592 13572 16596 13628
rect 16596 13572 16652 13628
rect 16652 13572 16656 13628
rect 16592 13568 16656 13572
rect 19352 13628 19416 13632
rect 19352 13572 19356 13628
rect 19356 13572 19412 13628
rect 19412 13572 19416 13628
rect 19352 13568 19416 13572
rect 19432 13628 19496 13632
rect 19432 13572 19436 13628
rect 19436 13572 19492 13628
rect 19492 13572 19496 13628
rect 19432 13568 19496 13572
rect 19512 13628 19576 13632
rect 19512 13572 19516 13628
rect 19516 13572 19572 13628
rect 19572 13572 19576 13628
rect 19512 13568 19576 13572
rect 19592 13628 19656 13632
rect 19592 13572 19596 13628
rect 19596 13572 19652 13628
rect 19652 13572 19656 13628
rect 19592 13568 19656 13572
rect 22352 13628 22416 13632
rect 22352 13572 22356 13628
rect 22356 13572 22412 13628
rect 22412 13572 22416 13628
rect 22352 13568 22416 13572
rect 22432 13628 22496 13632
rect 22432 13572 22436 13628
rect 22436 13572 22492 13628
rect 22492 13572 22496 13628
rect 22432 13568 22496 13572
rect 22512 13628 22576 13632
rect 22512 13572 22516 13628
rect 22516 13572 22572 13628
rect 22572 13572 22576 13628
rect 22512 13568 22576 13572
rect 22592 13628 22656 13632
rect 22592 13572 22596 13628
rect 22596 13572 22652 13628
rect 22652 13572 22656 13628
rect 22592 13568 22656 13572
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 2932 13084 2996 13088
rect 2932 13028 2936 13084
rect 2936 13028 2992 13084
rect 2992 13028 2996 13084
rect 2932 13024 2996 13028
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 5852 13084 5916 13088
rect 5852 13028 5856 13084
rect 5856 13028 5912 13084
rect 5912 13028 5916 13084
rect 5852 13024 5916 13028
rect 5932 13084 5996 13088
rect 5932 13028 5936 13084
rect 5936 13028 5992 13084
rect 5992 13028 5996 13084
rect 5932 13024 5996 13028
rect 6012 13084 6076 13088
rect 6012 13028 6016 13084
rect 6016 13028 6072 13084
rect 6072 13028 6076 13084
rect 6012 13024 6076 13028
rect 6092 13084 6156 13088
rect 6092 13028 6096 13084
rect 6096 13028 6152 13084
rect 6152 13028 6156 13084
rect 6092 13024 6156 13028
rect 8852 13084 8916 13088
rect 8852 13028 8856 13084
rect 8856 13028 8912 13084
rect 8912 13028 8916 13084
rect 8852 13024 8916 13028
rect 8932 13084 8996 13088
rect 8932 13028 8936 13084
rect 8936 13028 8992 13084
rect 8992 13028 8996 13084
rect 8932 13024 8996 13028
rect 9012 13084 9076 13088
rect 9012 13028 9016 13084
rect 9016 13028 9072 13084
rect 9072 13028 9076 13084
rect 9012 13024 9076 13028
rect 9092 13084 9156 13088
rect 9092 13028 9096 13084
rect 9096 13028 9152 13084
rect 9152 13028 9156 13084
rect 9092 13024 9156 13028
rect 11852 13084 11916 13088
rect 11852 13028 11856 13084
rect 11856 13028 11912 13084
rect 11912 13028 11916 13084
rect 11852 13024 11916 13028
rect 11932 13084 11996 13088
rect 11932 13028 11936 13084
rect 11936 13028 11992 13084
rect 11992 13028 11996 13084
rect 11932 13024 11996 13028
rect 12012 13084 12076 13088
rect 12012 13028 12016 13084
rect 12016 13028 12072 13084
rect 12072 13028 12076 13084
rect 12012 13024 12076 13028
rect 12092 13084 12156 13088
rect 12092 13028 12096 13084
rect 12096 13028 12152 13084
rect 12152 13028 12156 13084
rect 12092 13024 12156 13028
rect 14852 13084 14916 13088
rect 14852 13028 14856 13084
rect 14856 13028 14912 13084
rect 14912 13028 14916 13084
rect 14852 13024 14916 13028
rect 14932 13084 14996 13088
rect 14932 13028 14936 13084
rect 14936 13028 14992 13084
rect 14992 13028 14996 13084
rect 14932 13024 14996 13028
rect 15012 13084 15076 13088
rect 15012 13028 15016 13084
rect 15016 13028 15072 13084
rect 15072 13028 15076 13084
rect 15012 13024 15076 13028
rect 15092 13084 15156 13088
rect 15092 13028 15096 13084
rect 15096 13028 15152 13084
rect 15152 13028 15156 13084
rect 15092 13024 15156 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 17932 13084 17996 13088
rect 17932 13028 17936 13084
rect 17936 13028 17992 13084
rect 17992 13028 17996 13084
rect 17932 13024 17996 13028
rect 18012 13084 18076 13088
rect 18012 13028 18016 13084
rect 18016 13028 18072 13084
rect 18072 13028 18076 13084
rect 18012 13024 18076 13028
rect 18092 13084 18156 13088
rect 18092 13028 18096 13084
rect 18096 13028 18152 13084
rect 18152 13028 18156 13084
rect 18092 13024 18156 13028
rect 20852 13084 20916 13088
rect 20852 13028 20856 13084
rect 20856 13028 20912 13084
rect 20912 13028 20916 13084
rect 20852 13024 20916 13028
rect 20932 13084 20996 13088
rect 20932 13028 20936 13084
rect 20936 13028 20992 13084
rect 20992 13028 20996 13084
rect 20932 13024 20996 13028
rect 21012 13084 21076 13088
rect 21012 13028 21016 13084
rect 21016 13028 21072 13084
rect 21072 13028 21076 13084
rect 21012 13024 21076 13028
rect 21092 13084 21156 13088
rect 21092 13028 21096 13084
rect 21096 13028 21152 13084
rect 21152 13028 21156 13084
rect 21092 13024 21156 13028
rect 23852 13084 23916 13088
rect 23852 13028 23856 13084
rect 23856 13028 23912 13084
rect 23912 13028 23916 13084
rect 23852 13024 23916 13028
rect 23932 13084 23996 13088
rect 23932 13028 23936 13084
rect 23936 13028 23992 13084
rect 23992 13028 23996 13084
rect 23932 13024 23996 13028
rect 24012 13084 24076 13088
rect 24012 13028 24016 13084
rect 24016 13028 24072 13084
rect 24072 13028 24076 13084
rect 24012 13024 24076 13028
rect 24092 13084 24156 13088
rect 24092 13028 24096 13084
rect 24096 13028 24152 13084
rect 24152 13028 24156 13084
rect 24092 13024 24156 13028
rect 1352 12540 1416 12544
rect 1352 12484 1356 12540
rect 1356 12484 1412 12540
rect 1412 12484 1416 12540
rect 1352 12480 1416 12484
rect 1432 12540 1496 12544
rect 1432 12484 1436 12540
rect 1436 12484 1492 12540
rect 1492 12484 1496 12540
rect 1432 12480 1496 12484
rect 1512 12540 1576 12544
rect 1512 12484 1516 12540
rect 1516 12484 1572 12540
rect 1572 12484 1576 12540
rect 1512 12480 1576 12484
rect 1592 12540 1656 12544
rect 1592 12484 1596 12540
rect 1596 12484 1652 12540
rect 1652 12484 1656 12540
rect 1592 12480 1656 12484
rect 4352 12540 4416 12544
rect 4352 12484 4356 12540
rect 4356 12484 4412 12540
rect 4412 12484 4416 12540
rect 4352 12480 4416 12484
rect 4432 12540 4496 12544
rect 4432 12484 4436 12540
rect 4436 12484 4492 12540
rect 4492 12484 4496 12540
rect 4432 12480 4496 12484
rect 4512 12540 4576 12544
rect 4512 12484 4516 12540
rect 4516 12484 4572 12540
rect 4572 12484 4576 12540
rect 4512 12480 4576 12484
rect 4592 12540 4656 12544
rect 4592 12484 4596 12540
rect 4596 12484 4652 12540
rect 4652 12484 4656 12540
rect 4592 12480 4656 12484
rect 7352 12540 7416 12544
rect 7352 12484 7356 12540
rect 7356 12484 7412 12540
rect 7412 12484 7416 12540
rect 7352 12480 7416 12484
rect 7432 12540 7496 12544
rect 7432 12484 7436 12540
rect 7436 12484 7492 12540
rect 7492 12484 7496 12540
rect 7432 12480 7496 12484
rect 7512 12540 7576 12544
rect 7512 12484 7516 12540
rect 7516 12484 7572 12540
rect 7572 12484 7576 12540
rect 7512 12480 7576 12484
rect 7592 12540 7656 12544
rect 7592 12484 7596 12540
rect 7596 12484 7652 12540
rect 7652 12484 7656 12540
rect 7592 12480 7656 12484
rect 10352 12540 10416 12544
rect 10352 12484 10356 12540
rect 10356 12484 10412 12540
rect 10412 12484 10416 12540
rect 10352 12480 10416 12484
rect 10432 12540 10496 12544
rect 10432 12484 10436 12540
rect 10436 12484 10492 12540
rect 10492 12484 10496 12540
rect 10432 12480 10496 12484
rect 10512 12540 10576 12544
rect 10512 12484 10516 12540
rect 10516 12484 10572 12540
rect 10572 12484 10576 12540
rect 10512 12480 10576 12484
rect 10592 12540 10656 12544
rect 10592 12484 10596 12540
rect 10596 12484 10652 12540
rect 10652 12484 10656 12540
rect 10592 12480 10656 12484
rect 13352 12540 13416 12544
rect 13352 12484 13356 12540
rect 13356 12484 13412 12540
rect 13412 12484 13416 12540
rect 13352 12480 13416 12484
rect 13432 12540 13496 12544
rect 13432 12484 13436 12540
rect 13436 12484 13492 12540
rect 13492 12484 13496 12540
rect 13432 12480 13496 12484
rect 13512 12540 13576 12544
rect 13512 12484 13516 12540
rect 13516 12484 13572 12540
rect 13572 12484 13576 12540
rect 13512 12480 13576 12484
rect 13592 12540 13656 12544
rect 13592 12484 13596 12540
rect 13596 12484 13652 12540
rect 13652 12484 13656 12540
rect 13592 12480 13656 12484
rect 16352 12540 16416 12544
rect 16352 12484 16356 12540
rect 16356 12484 16412 12540
rect 16412 12484 16416 12540
rect 16352 12480 16416 12484
rect 16432 12540 16496 12544
rect 16432 12484 16436 12540
rect 16436 12484 16492 12540
rect 16492 12484 16496 12540
rect 16432 12480 16496 12484
rect 16512 12540 16576 12544
rect 16512 12484 16516 12540
rect 16516 12484 16572 12540
rect 16572 12484 16576 12540
rect 16512 12480 16576 12484
rect 16592 12540 16656 12544
rect 16592 12484 16596 12540
rect 16596 12484 16652 12540
rect 16652 12484 16656 12540
rect 16592 12480 16656 12484
rect 19352 12540 19416 12544
rect 19352 12484 19356 12540
rect 19356 12484 19412 12540
rect 19412 12484 19416 12540
rect 19352 12480 19416 12484
rect 19432 12540 19496 12544
rect 19432 12484 19436 12540
rect 19436 12484 19492 12540
rect 19492 12484 19496 12540
rect 19432 12480 19496 12484
rect 19512 12540 19576 12544
rect 19512 12484 19516 12540
rect 19516 12484 19572 12540
rect 19572 12484 19576 12540
rect 19512 12480 19576 12484
rect 19592 12540 19656 12544
rect 19592 12484 19596 12540
rect 19596 12484 19652 12540
rect 19652 12484 19656 12540
rect 19592 12480 19656 12484
rect 22352 12540 22416 12544
rect 22352 12484 22356 12540
rect 22356 12484 22412 12540
rect 22412 12484 22416 12540
rect 22352 12480 22416 12484
rect 22432 12540 22496 12544
rect 22432 12484 22436 12540
rect 22436 12484 22492 12540
rect 22492 12484 22496 12540
rect 22432 12480 22496 12484
rect 22512 12540 22576 12544
rect 22512 12484 22516 12540
rect 22516 12484 22572 12540
rect 22572 12484 22576 12540
rect 22512 12480 22576 12484
rect 22592 12540 22656 12544
rect 22592 12484 22596 12540
rect 22596 12484 22652 12540
rect 22652 12484 22656 12540
rect 22592 12480 22656 12484
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 2932 11996 2996 12000
rect 2932 11940 2936 11996
rect 2936 11940 2992 11996
rect 2992 11940 2996 11996
rect 2932 11936 2996 11940
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 5852 11996 5916 12000
rect 5852 11940 5856 11996
rect 5856 11940 5912 11996
rect 5912 11940 5916 11996
rect 5852 11936 5916 11940
rect 5932 11996 5996 12000
rect 5932 11940 5936 11996
rect 5936 11940 5992 11996
rect 5992 11940 5996 11996
rect 5932 11936 5996 11940
rect 6012 11996 6076 12000
rect 6012 11940 6016 11996
rect 6016 11940 6072 11996
rect 6072 11940 6076 11996
rect 6012 11936 6076 11940
rect 6092 11996 6156 12000
rect 6092 11940 6096 11996
rect 6096 11940 6152 11996
rect 6152 11940 6156 11996
rect 6092 11936 6156 11940
rect 8852 11996 8916 12000
rect 8852 11940 8856 11996
rect 8856 11940 8912 11996
rect 8912 11940 8916 11996
rect 8852 11936 8916 11940
rect 8932 11996 8996 12000
rect 8932 11940 8936 11996
rect 8936 11940 8992 11996
rect 8992 11940 8996 11996
rect 8932 11936 8996 11940
rect 9012 11996 9076 12000
rect 9012 11940 9016 11996
rect 9016 11940 9072 11996
rect 9072 11940 9076 11996
rect 9012 11936 9076 11940
rect 9092 11996 9156 12000
rect 9092 11940 9096 11996
rect 9096 11940 9152 11996
rect 9152 11940 9156 11996
rect 9092 11936 9156 11940
rect 11852 11996 11916 12000
rect 11852 11940 11856 11996
rect 11856 11940 11912 11996
rect 11912 11940 11916 11996
rect 11852 11936 11916 11940
rect 11932 11996 11996 12000
rect 11932 11940 11936 11996
rect 11936 11940 11992 11996
rect 11992 11940 11996 11996
rect 11932 11936 11996 11940
rect 12012 11996 12076 12000
rect 12012 11940 12016 11996
rect 12016 11940 12072 11996
rect 12072 11940 12076 11996
rect 12012 11936 12076 11940
rect 12092 11996 12156 12000
rect 12092 11940 12096 11996
rect 12096 11940 12152 11996
rect 12152 11940 12156 11996
rect 12092 11936 12156 11940
rect 14852 11996 14916 12000
rect 14852 11940 14856 11996
rect 14856 11940 14912 11996
rect 14912 11940 14916 11996
rect 14852 11936 14916 11940
rect 14932 11996 14996 12000
rect 14932 11940 14936 11996
rect 14936 11940 14992 11996
rect 14992 11940 14996 11996
rect 14932 11936 14996 11940
rect 15012 11996 15076 12000
rect 15012 11940 15016 11996
rect 15016 11940 15072 11996
rect 15072 11940 15076 11996
rect 15012 11936 15076 11940
rect 15092 11996 15156 12000
rect 15092 11940 15096 11996
rect 15096 11940 15152 11996
rect 15152 11940 15156 11996
rect 15092 11936 15156 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 17932 11996 17996 12000
rect 17932 11940 17936 11996
rect 17936 11940 17992 11996
rect 17992 11940 17996 11996
rect 17932 11936 17996 11940
rect 18012 11996 18076 12000
rect 18012 11940 18016 11996
rect 18016 11940 18072 11996
rect 18072 11940 18076 11996
rect 18012 11936 18076 11940
rect 18092 11996 18156 12000
rect 18092 11940 18096 11996
rect 18096 11940 18152 11996
rect 18152 11940 18156 11996
rect 18092 11936 18156 11940
rect 20852 11996 20916 12000
rect 20852 11940 20856 11996
rect 20856 11940 20912 11996
rect 20912 11940 20916 11996
rect 20852 11936 20916 11940
rect 20932 11996 20996 12000
rect 20932 11940 20936 11996
rect 20936 11940 20992 11996
rect 20992 11940 20996 11996
rect 20932 11936 20996 11940
rect 21012 11996 21076 12000
rect 21012 11940 21016 11996
rect 21016 11940 21072 11996
rect 21072 11940 21076 11996
rect 21012 11936 21076 11940
rect 21092 11996 21156 12000
rect 21092 11940 21096 11996
rect 21096 11940 21152 11996
rect 21152 11940 21156 11996
rect 21092 11936 21156 11940
rect 23852 11996 23916 12000
rect 23852 11940 23856 11996
rect 23856 11940 23912 11996
rect 23912 11940 23916 11996
rect 23852 11936 23916 11940
rect 23932 11996 23996 12000
rect 23932 11940 23936 11996
rect 23936 11940 23992 11996
rect 23992 11940 23996 11996
rect 23932 11936 23996 11940
rect 24012 11996 24076 12000
rect 24012 11940 24016 11996
rect 24016 11940 24072 11996
rect 24072 11940 24076 11996
rect 24012 11936 24076 11940
rect 24092 11996 24156 12000
rect 24092 11940 24096 11996
rect 24096 11940 24152 11996
rect 24152 11940 24156 11996
rect 24092 11936 24156 11940
rect 1352 11452 1416 11456
rect 1352 11396 1356 11452
rect 1356 11396 1412 11452
rect 1412 11396 1416 11452
rect 1352 11392 1416 11396
rect 1432 11452 1496 11456
rect 1432 11396 1436 11452
rect 1436 11396 1492 11452
rect 1492 11396 1496 11452
rect 1432 11392 1496 11396
rect 1512 11452 1576 11456
rect 1512 11396 1516 11452
rect 1516 11396 1572 11452
rect 1572 11396 1576 11452
rect 1512 11392 1576 11396
rect 1592 11452 1656 11456
rect 1592 11396 1596 11452
rect 1596 11396 1652 11452
rect 1652 11396 1656 11452
rect 1592 11392 1656 11396
rect 4352 11452 4416 11456
rect 4352 11396 4356 11452
rect 4356 11396 4412 11452
rect 4412 11396 4416 11452
rect 4352 11392 4416 11396
rect 4432 11452 4496 11456
rect 4432 11396 4436 11452
rect 4436 11396 4492 11452
rect 4492 11396 4496 11452
rect 4432 11392 4496 11396
rect 4512 11452 4576 11456
rect 4512 11396 4516 11452
rect 4516 11396 4572 11452
rect 4572 11396 4576 11452
rect 4512 11392 4576 11396
rect 4592 11452 4656 11456
rect 4592 11396 4596 11452
rect 4596 11396 4652 11452
rect 4652 11396 4656 11452
rect 4592 11392 4656 11396
rect 7352 11452 7416 11456
rect 7352 11396 7356 11452
rect 7356 11396 7412 11452
rect 7412 11396 7416 11452
rect 7352 11392 7416 11396
rect 7432 11452 7496 11456
rect 7432 11396 7436 11452
rect 7436 11396 7492 11452
rect 7492 11396 7496 11452
rect 7432 11392 7496 11396
rect 7512 11452 7576 11456
rect 7512 11396 7516 11452
rect 7516 11396 7572 11452
rect 7572 11396 7576 11452
rect 7512 11392 7576 11396
rect 7592 11452 7656 11456
rect 7592 11396 7596 11452
rect 7596 11396 7652 11452
rect 7652 11396 7656 11452
rect 7592 11392 7656 11396
rect 10352 11452 10416 11456
rect 10352 11396 10356 11452
rect 10356 11396 10412 11452
rect 10412 11396 10416 11452
rect 10352 11392 10416 11396
rect 10432 11452 10496 11456
rect 10432 11396 10436 11452
rect 10436 11396 10492 11452
rect 10492 11396 10496 11452
rect 10432 11392 10496 11396
rect 10512 11452 10576 11456
rect 10512 11396 10516 11452
rect 10516 11396 10572 11452
rect 10572 11396 10576 11452
rect 10512 11392 10576 11396
rect 10592 11452 10656 11456
rect 10592 11396 10596 11452
rect 10596 11396 10652 11452
rect 10652 11396 10656 11452
rect 10592 11392 10656 11396
rect 13352 11452 13416 11456
rect 13352 11396 13356 11452
rect 13356 11396 13412 11452
rect 13412 11396 13416 11452
rect 13352 11392 13416 11396
rect 13432 11452 13496 11456
rect 13432 11396 13436 11452
rect 13436 11396 13492 11452
rect 13492 11396 13496 11452
rect 13432 11392 13496 11396
rect 13512 11452 13576 11456
rect 13512 11396 13516 11452
rect 13516 11396 13572 11452
rect 13572 11396 13576 11452
rect 13512 11392 13576 11396
rect 13592 11452 13656 11456
rect 13592 11396 13596 11452
rect 13596 11396 13652 11452
rect 13652 11396 13656 11452
rect 13592 11392 13656 11396
rect 16352 11452 16416 11456
rect 16352 11396 16356 11452
rect 16356 11396 16412 11452
rect 16412 11396 16416 11452
rect 16352 11392 16416 11396
rect 16432 11452 16496 11456
rect 16432 11396 16436 11452
rect 16436 11396 16492 11452
rect 16492 11396 16496 11452
rect 16432 11392 16496 11396
rect 16512 11452 16576 11456
rect 16512 11396 16516 11452
rect 16516 11396 16572 11452
rect 16572 11396 16576 11452
rect 16512 11392 16576 11396
rect 16592 11452 16656 11456
rect 16592 11396 16596 11452
rect 16596 11396 16652 11452
rect 16652 11396 16656 11452
rect 16592 11392 16656 11396
rect 19352 11452 19416 11456
rect 19352 11396 19356 11452
rect 19356 11396 19412 11452
rect 19412 11396 19416 11452
rect 19352 11392 19416 11396
rect 19432 11452 19496 11456
rect 19432 11396 19436 11452
rect 19436 11396 19492 11452
rect 19492 11396 19496 11452
rect 19432 11392 19496 11396
rect 19512 11452 19576 11456
rect 19512 11396 19516 11452
rect 19516 11396 19572 11452
rect 19572 11396 19576 11452
rect 19512 11392 19576 11396
rect 19592 11452 19656 11456
rect 19592 11396 19596 11452
rect 19596 11396 19652 11452
rect 19652 11396 19656 11452
rect 19592 11392 19656 11396
rect 22352 11452 22416 11456
rect 22352 11396 22356 11452
rect 22356 11396 22412 11452
rect 22412 11396 22416 11452
rect 22352 11392 22416 11396
rect 22432 11452 22496 11456
rect 22432 11396 22436 11452
rect 22436 11396 22492 11452
rect 22492 11396 22496 11452
rect 22432 11392 22496 11396
rect 22512 11452 22576 11456
rect 22512 11396 22516 11452
rect 22516 11396 22572 11452
rect 22572 11396 22576 11452
rect 22512 11392 22576 11396
rect 22592 11452 22656 11456
rect 22592 11396 22596 11452
rect 22596 11396 22652 11452
rect 22652 11396 22656 11452
rect 22592 11392 22656 11396
rect 13124 11052 13188 11116
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 2932 10908 2996 10912
rect 2932 10852 2936 10908
rect 2936 10852 2992 10908
rect 2992 10852 2996 10908
rect 2932 10848 2996 10852
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 5852 10908 5916 10912
rect 5852 10852 5856 10908
rect 5856 10852 5912 10908
rect 5912 10852 5916 10908
rect 5852 10848 5916 10852
rect 5932 10908 5996 10912
rect 5932 10852 5936 10908
rect 5936 10852 5992 10908
rect 5992 10852 5996 10908
rect 5932 10848 5996 10852
rect 6012 10908 6076 10912
rect 6012 10852 6016 10908
rect 6016 10852 6072 10908
rect 6072 10852 6076 10908
rect 6012 10848 6076 10852
rect 6092 10908 6156 10912
rect 6092 10852 6096 10908
rect 6096 10852 6152 10908
rect 6152 10852 6156 10908
rect 6092 10848 6156 10852
rect 8852 10908 8916 10912
rect 8852 10852 8856 10908
rect 8856 10852 8912 10908
rect 8912 10852 8916 10908
rect 8852 10848 8916 10852
rect 8932 10908 8996 10912
rect 8932 10852 8936 10908
rect 8936 10852 8992 10908
rect 8992 10852 8996 10908
rect 8932 10848 8996 10852
rect 9012 10908 9076 10912
rect 9012 10852 9016 10908
rect 9016 10852 9072 10908
rect 9072 10852 9076 10908
rect 9012 10848 9076 10852
rect 9092 10908 9156 10912
rect 9092 10852 9096 10908
rect 9096 10852 9152 10908
rect 9152 10852 9156 10908
rect 9092 10848 9156 10852
rect 11852 10908 11916 10912
rect 11852 10852 11856 10908
rect 11856 10852 11912 10908
rect 11912 10852 11916 10908
rect 11852 10848 11916 10852
rect 11932 10908 11996 10912
rect 11932 10852 11936 10908
rect 11936 10852 11992 10908
rect 11992 10852 11996 10908
rect 11932 10848 11996 10852
rect 12012 10908 12076 10912
rect 12012 10852 12016 10908
rect 12016 10852 12072 10908
rect 12072 10852 12076 10908
rect 12012 10848 12076 10852
rect 12092 10908 12156 10912
rect 12092 10852 12096 10908
rect 12096 10852 12152 10908
rect 12152 10852 12156 10908
rect 12092 10848 12156 10852
rect 14852 10908 14916 10912
rect 14852 10852 14856 10908
rect 14856 10852 14912 10908
rect 14912 10852 14916 10908
rect 14852 10848 14916 10852
rect 14932 10908 14996 10912
rect 14932 10852 14936 10908
rect 14936 10852 14992 10908
rect 14992 10852 14996 10908
rect 14932 10848 14996 10852
rect 15012 10908 15076 10912
rect 15012 10852 15016 10908
rect 15016 10852 15072 10908
rect 15072 10852 15076 10908
rect 15012 10848 15076 10852
rect 15092 10908 15156 10912
rect 15092 10852 15096 10908
rect 15096 10852 15152 10908
rect 15152 10852 15156 10908
rect 15092 10848 15156 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 17932 10908 17996 10912
rect 17932 10852 17936 10908
rect 17936 10852 17992 10908
rect 17992 10852 17996 10908
rect 17932 10848 17996 10852
rect 18012 10908 18076 10912
rect 18012 10852 18016 10908
rect 18016 10852 18072 10908
rect 18072 10852 18076 10908
rect 18012 10848 18076 10852
rect 18092 10908 18156 10912
rect 18092 10852 18096 10908
rect 18096 10852 18152 10908
rect 18152 10852 18156 10908
rect 18092 10848 18156 10852
rect 20852 10908 20916 10912
rect 20852 10852 20856 10908
rect 20856 10852 20912 10908
rect 20912 10852 20916 10908
rect 20852 10848 20916 10852
rect 20932 10908 20996 10912
rect 20932 10852 20936 10908
rect 20936 10852 20992 10908
rect 20992 10852 20996 10908
rect 20932 10848 20996 10852
rect 21012 10908 21076 10912
rect 21012 10852 21016 10908
rect 21016 10852 21072 10908
rect 21072 10852 21076 10908
rect 21012 10848 21076 10852
rect 21092 10908 21156 10912
rect 21092 10852 21096 10908
rect 21096 10852 21152 10908
rect 21152 10852 21156 10908
rect 21092 10848 21156 10852
rect 23852 10908 23916 10912
rect 23852 10852 23856 10908
rect 23856 10852 23912 10908
rect 23912 10852 23916 10908
rect 23852 10848 23916 10852
rect 23932 10908 23996 10912
rect 23932 10852 23936 10908
rect 23936 10852 23992 10908
rect 23992 10852 23996 10908
rect 23932 10848 23996 10852
rect 24012 10908 24076 10912
rect 24012 10852 24016 10908
rect 24016 10852 24072 10908
rect 24072 10852 24076 10908
rect 24012 10848 24076 10852
rect 24092 10908 24156 10912
rect 24092 10852 24096 10908
rect 24096 10852 24152 10908
rect 24152 10852 24156 10908
rect 24092 10848 24156 10852
rect 1352 10364 1416 10368
rect 1352 10308 1356 10364
rect 1356 10308 1412 10364
rect 1412 10308 1416 10364
rect 1352 10304 1416 10308
rect 1432 10364 1496 10368
rect 1432 10308 1436 10364
rect 1436 10308 1492 10364
rect 1492 10308 1496 10364
rect 1432 10304 1496 10308
rect 1512 10364 1576 10368
rect 1512 10308 1516 10364
rect 1516 10308 1572 10364
rect 1572 10308 1576 10364
rect 1512 10304 1576 10308
rect 1592 10364 1656 10368
rect 1592 10308 1596 10364
rect 1596 10308 1652 10364
rect 1652 10308 1656 10364
rect 1592 10304 1656 10308
rect 4352 10364 4416 10368
rect 4352 10308 4356 10364
rect 4356 10308 4412 10364
rect 4412 10308 4416 10364
rect 4352 10304 4416 10308
rect 4432 10364 4496 10368
rect 4432 10308 4436 10364
rect 4436 10308 4492 10364
rect 4492 10308 4496 10364
rect 4432 10304 4496 10308
rect 4512 10364 4576 10368
rect 4512 10308 4516 10364
rect 4516 10308 4572 10364
rect 4572 10308 4576 10364
rect 4512 10304 4576 10308
rect 4592 10364 4656 10368
rect 4592 10308 4596 10364
rect 4596 10308 4652 10364
rect 4652 10308 4656 10364
rect 4592 10304 4656 10308
rect 7352 10364 7416 10368
rect 7352 10308 7356 10364
rect 7356 10308 7412 10364
rect 7412 10308 7416 10364
rect 7352 10304 7416 10308
rect 7432 10364 7496 10368
rect 7432 10308 7436 10364
rect 7436 10308 7492 10364
rect 7492 10308 7496 10364
rect 7432 10304 7496 10308
rect 7512 10364 7576 10368
rect 7512 10308 7516 10364
rect 7516 10308 7572 10364
rect 7572 10308 7576 10364
rect 7512 10304 7576 10308
rect 7592 10364 7656 10368
rect 7592 10308 7596 10364
rect 7596 10308 7652 10364
rect 7652 10308 7656 10364
rect 7592 10304 7656 10308
rect 10352 10364 10416 10368
rect 10352 10308 10356 10364
rect 10356 10308 10412 10364
rect 10412 10308 10416 10364
rect 10352 10304 10416 10308
rect 10432 10364 10496 10368
rect 10432 10308 10436 10364
rect 10436 10308 10492 10364
rect 10492 10308 10496 10364
rect 10432 10304 10496 10308
rect 10512 10364 10576 10368
rect 10512 10308 10516 10364
rect 10516 10308 10572 10364
rect 10572 10308 10576 10364
rect 10512 10304 10576 10308
rect 10592 10364 10656 10368
rect 10592 10308 10596 10364
rect 10596 10308 10652 10364
rect 10652 10308 10656 10364
rect 10592 10304 10656 10308
rect 13352 10364 13416 10368
rect 13352 10308 13356 10364
rect 13356 10308 13412 10364
rect 13412 10308 13416 10364
rect 13352 10304 13416 10308
rect 13432 10364 13496 10368
rect 13432 10308 13436 10364
rect 13436 10308 13492 10364
rect 13492 10308 13496 10364
rect 13432 10304 13496 10308
rect 13512 10364 13576 10368
rect 13512 10308 13516 10364
rect 13516 10308 13572 10364
rect 13572 10308 13576 10364
rect 13512 10304 13576 10308
rect 13592 10364 13656 10368
rect 13592 10308 13596 10364
rect 13596 10308 13652 10364
rect 13652 10308 13656 10364
rect 13592 10304 13656 10308
rect 16352 10364 16416 10368
rect 16352 10308 16356 10364
rect 16356 10308 16412 10364
rect 16412 10308 16416 10364
rect 16352 10304 16416 10308
rect 16432 10364 16496 10368
rect 16432 10308 16436 10364
rect 16436 10308 16492 10364
rect 16492 10308 16496 10364
rect 16432 10304 16496 10308
rect 16512 10364 16576 10368
rect 16512 10308 16516 10364
rect 16516 10308 16572 10364
rect 16572 10308 16576 10364
rect 16512 10304 16576 10308
rect 16592 10364 16656 10368
rect 16592 10308 16596 10364
rect 16596 10308 16652 10364
rect 16652 10308 16656 10364
rect 16592 10304 16656 10308
rect 19352 10364 19416 10368
rect 19352 10308 19356 10364
rect 19356 10308 19412 10364
rect 19412 10308 19416 10364
rect 19352 10304 19416 10308
rect 19432 10364 19496 10368
rect 19432 10308 19436 10364
rect 19436 10308 19492 10364
rect 19492 10308 19496 10364
rect 19432 10304 19496 10308
rect 19512 10364 19576 10368
rect 19512 10308 19516 10364
rect 19516 10308 19572 10364
rect 19572 10308 19576 10364
rect 19512 10304 19576 10308
rect 19592 10364 19656 10368
rect 19592 10308 19596 10364
rect 19596 10308 19652 10364
rect 19652 10308 19656 10364
rect 19592 10304 19656 10308
rect 22352 10364 22416 10368
rect 22352 10308 22356 10364
rect 22356 10308 22412 10364
rect 22412 10308 22416 10364
rect 22352 10304 22416 10308
rect 22432 10364 22496 10368
rect 22432 10308 22436 10364
rect 22436 10308 22492 10364
rect 22492 10308 22496 10364
rect 22432 10304 22496 10308
rect 22512 10364 22576 10368
rect 22512 10308 22516 10364
rect 22516 10308 22572 10364
rect 22572 10308 22576 10364
rect 22512 10304 22576 10308
rect 22592 10364 22656 10368
rect 22592 10308 22596 10364
rect 22596 10308 22652 10364
rect 22652 10308 22656 10364
rect 22592 10304 22656 10308
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 2932 9820 2996 9824
rect 2932 9764 2936 9820
rect 2936 9764 2992 9820
rect 2992 9764 2996 9820
rect 2932 9760 2996 9764
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 5852 9820 5916 9824
rect 5852 9764 5856 9820
rect 5856 9764 5912 9820
rect 5912 9764 5916 9820
rect 5852 9760 5916 9764
rect 5932 9820 5996 9824
rect 5932 9764 5936 9820
rect 5936 9764 5992 9820
rect 5992 9764 5996 9820
rect 5932 9760 5996 9764
rect 6012 9820 6076 9824
rect 6012 9764 6016 9820
rect 6016 9764 6072 9820
rect 6072 9764 6076 9820
rect 6012 9760 6076 9764
rect 6092 9820 6156 9824
rect 6092 9764 6096 9820
rect 6096 9764 6152 9820
rect 6152 9764 6156 9820
rect 6092 9760 6156 9764
rect 8852 9820 8916 9824
rect 8852 9764 8856 9820
rect 8856 9764 8912 9820
rect 8912 9764 8916 9820
rect 8852 9760 8916 9764
rect 8932 9820 8996 9824
rect 8932 9764 8936 9820
rect 8936 9764 8992 9820
rect 8992 9764 8996 9820
rect 8932 9760 8996 9764
rect 9012 9820 9076 9824
rect 9012 9764 9016 9820
rect 9016 9764 9072 9820
rect 9072 9764 9076 9820
rect 9012 9760 9076 9764
rect 9092 9820 9156 9824
rect 9092 9764 9096 9820
rect 9096 9764 9152 9820
rect 9152 9764 9156 9820
rect 9092 9760 9156 9764
rect 11852 9820 11916 9824
rect 11852 9764 11856 9820
rect 11856 9764 11912 9820
rect 11912 9764 11916 9820
rect 11852 9760 11916 9764
rect 11932 9820 11996 9824
rect 11932 9764 11936 9820
rect 11936 9764 11992 9820
rect 11992 9764 11996 9820
rect 11932 9760 11996 9764
rect 12012 9820 12076 9824
rect 12012 9764 12016 9820
rect 12016 9764 12072 9820
rect 12072 9764 12076 9820
rect 12012 9760 12076 9764
rect 12092 9820 12156 9824
rect 12092 9764 12096 9820
rect 12096 9764 12152 9820
rect 12152 9764 12156 9820
rect 12092 9760 12156 9764
rect 14852 9820 14916 9824
rect 14852 9764 14856 9820
rect 14856 9764 14912 9820
rect 14912 9764 14916 9820
rect 14852 9760 14916 9764
rect 14932 9820 14996 9824
rect 14932 9764 14936 9820
rect 14936 9764 14992 9820
rect 14992 9764 14996 9820
rect 14932 9760 14996 9764
rect 15012 9820 15076 9824
rect 15012 9764 15016 9820
rect 15016 9764 15072 9820
rect 15072 9764 15076 9820
rect 15012 9760 15076 9764
rect 15092 9820 15156 9824
rect 15092 9764 15096 9820
rect 15096 9764 15152 9820
rect 15152 9764 15156 9820
rect 15092 9760 15156 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 17932 9820 17996 9824
rect 17932 9764 17936 9820
rect 17936 9764 17992 9820
rect 17992 9764 17996 9820
rect 17932 9760 17996 9764
rect 18012 9820 18076 9824
rect 18012 9764 18016 9820
rect 18016 9764 18072 9820
rect 18072 9764 18076 9820
rect 18012 9760 18076 9764
rect 18092 9820 18156 9824
rect 18092 9764 18096 9820
rect 18096 9764 18152 9820
rect 18152 9764 18156 9820
rect 18092 9760 18156 9764
rect 20852 9820 20916 9824
rect 20852 9764 20856 9820
rect 20856 9764 20912 9820
rect 20912 9764 20916 9820
rect 20852 9760 20916 9764
rect 20932 9820 20996 9824
rect 20932 9764 20936 9820
rect 20936 9764 20992 9820
rect 20992 9764 20996 9820
rect 20932 9760 20996 9764
rect 21012 9820 21076 9824
rect 21012 9764 21016 9820
rect 21016 9764 21072 9820
rect 21072 9764 21076 9820
rect 21012 9760 21076 9764
rect 21092 9820 21156 9824
rect 21092 9764 21096 9820
rect 21096 9764 21152 9820
rect 21152 9764 21156 9820
rect 21092 9760 21156 9764
rect 23852 9820 23916 9824
rect 23852 9764 23856 9820
rect 23856 9764 23912 9820
rect 23912 9764 23916 9820
rect 23852 9760 23916 9764
rect 23932 9820 23996 9824
rect 23932 9764 23936 9820
rect 23936 9764 23992 9820
rect 23992 9764 23996 9820
rect 23932 9760 23996 9764
rect 24012 9820 24076 9824
rect 24012 9764 24016 9820
rect 24016 9764 24072 9820
rect 24072 9764 24076 9820
rect 24012 9760 24076 9764
rect 24092 9820 24156 9824
rect 24092 9764 24096 9820
rect 24096 9764 24152 9820
rect 24152 9764 24156 9820
rect 24092 9760 24156 9764
rect 1352 9276 1416 9280
rect 1352 9220 1356 9276
rect 1356 9220 1412 9276
rect 1412 9220 1416 9276
rect 1352 9216 1416 9220
rect 1432 9276 1496 9280
rect 1432 9220 1436 9276
rect 1436 9220 1492 9276
rect 1492 9220 1496 9276
rect 1432 9216 1496 9220
rect 1512 9276 1576 9280
rect 1512 9220 1516 9276
rect 1516 9220 1572 9276
rect 1572 9220 1576 9276
rect 1512 9216 1576 9220
rect 1592 9276 1656 9280
rect 1592 9220 1596 9276
rect 1596 9220 1652 9276
rect 1652 9220 1656 9276
rect 1592 9216 1656 9220
rect 4352 9276 4416 9280
rect 4352 9220 4356 9276
rect 4356 9220 4412 9276
rect 4412 9220 4416 9276
rect 4352 9216 4416 9220
rect 4432 9276 4496 9280
rect 4432 9220 4436 9276
rect 4436 9220 4492 9276
rect 4492 9220 4496 9276
rect 4432 9216 4496 9220
rect 4512 9276 4576 9280
rect 4512 9220 4516 9276
rect 4516 9220 4572 9276
rect 4572 9220 4576 9276
rect 4512 9216 4576 9220
rect 4592 9276 4656 9280
rect 4592 9220 4596 9276
rect 4596 9220 4652 9276
rect 4652 9220 4656 9276
rect 4592 9216 4656 9220
rect 7352 9276 7416 9280
rect 7352 9220 7356 9276
rect 7356 9220 7412 9276
rect 7412 9220 7416 9276
rect 7352 9216 7416 9220
rect 7432 9276 7496 9280
rect 7432 9220 7436 9276
rect 7436 9220 7492 9276
rect 7492 9220 7496 9276
rect 7432 9216 7496 9220
rect 7512 9276 7576 9280
rect 7512 9220 7516 9276
rect 7516 9220 7572 9276
rect 7572 9220 7576 9276
rect 7512 9216 7576 9220
rect 7592 9276 7656 9280
rect 7592 9220 7596 9276
rect 7596 9220 7652 9276
rect 7652 9220 7656 9276
rect 7592 9216 7656 9220
rect 10352 9276 10416 9280
rect 10352 9220 10356 9276
rect 10356 9220 10412 9276
rect 10412 9220 10416 9276
rect 10352 9216 10416 9220
rect 10432 9276 10496 9280
rect 10432 9220 10436 9276
rect 10436 9220 10492 9276
rect 10492 9220 10496 9276
rect 10432 9216 10496 9220
rect 10512 9276 10576 9280
rect 10512 9220 10516 9276
rect 10516 9220 10572 9276
rect 10572 9220 10576 9276
rect 10512 9216 10576 9220
rect 10592 9276 10656 9280
rect 10592 9220 10596 9276
rect 10596 9220 10652 9276
rect 10652 9220 10656 9276
rect 10592 9216 10656 9220
rect 13352 9276 13416 9280
rect 13352 9220 13356 9276
rect 13356 9220 13412 9276
rect 13412 9220 13416 9276
rect 13352 9216 13416 9220
rect 13432 9276 13496 9280
rect 13432 9220 13436 9276
rect 13436 9220 13492 9276
rect 13492 9220 13496 9276
rect 13432 9216 13496 9220
rect 13512 9276 13576 9280
rect 13512 9220 13516 9276
rect 13516 9220 13572 9276
rect 13572 9220 13576 9276
rect 13512 9216 13576 9220
rect 13592 9276 13656 9280
rect 13592 9220 13596 9276
rect 13596 9220 13652 9276
rect 13652 9220 13656 9276
rect 13592 9216 13656 9220
rect 16352 9276 16416 9280
rect 16352 9220 16356 9276
rect 16356 9220 16412 9276
rect 16412 9220 16416 9276
rect 16352 9216 16416 9220
rect 16432 9276 16496 9280
rect 16432 9220 16436 9276
rect 16436 9220 16492 9276
rect 16492 9220 16496 9276
rect 16432 9216 16496 9220
rect 16512 9276 16576 9280
rect 16512 9220 16516 9276
rect 16516 9220 16572 9276
rect 16572 9220 16576 9276
rect 16512 9216 16576 9220
rect 16592 9276 16656 9280
rect 16592 9220 16596 9276
rect 16596 9220 16652 9276
rect 16652 9220 16656 9276
rect 16592 9216 16656 9220
rect 19352 9276 19416 9280
rect 19352 9220 19356 9276
rect 19356 9220 19412 9276
rect 19412 9220 19416 9276
rect 19352 9216 19416 9220
rect 19432 9276 19496 9280
rect 19432 9220 19436 9276
rect 19436 9220 19492 9276
rect 19492 9220 19496 9276
rect 19432 9216 19496 9220
rect 19512 9276 19576 9280
rect 19512 9220 19516 9276
rect 19516 9220 19572 9276
rect 19572 9220 19576 9276
rect 19512 9216 19576 9220
rect 19592 9276 19656 9280
rect 19592 9220 19596 9276
rect 19596 9220 19652 9276
rect 19652 9220 19656 9276
rect 19592 9216 19656 9220
rect 22352 9276 22416 9280
rect 22352 9220 22356 9276
rect 22356 9220 22412 9276
rect 22412 9220 22416 9276
rect 22352 9216 22416 9220
rect 22432 9276 22496 9280
rect 22432 9220 22436 9276
rect 22436 9220 22492 9276
rect 22492 9220 22496 9276
rect 22432 9216 22496 9220
rect 22512 9276 22576 9280
rect 22512 9220 22516 9276
rect 22516 9220 22572 9276
rect 22572 9220 22576 9276
rect 22512 9216 22576 9220
rect 22592 9276 22656 9280
rect 22592 9220 22596 9276
rect 22596 9220 22652 9276
rect 22652 9220 22656 9276
rect 22592 9216 22656 9220
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 2932 8732 2996 8736
rect 2932 8676 2936 8732
rect 2936 8676 2992 8732
rect 2992 8676 2996 8732
rect 2932 8672 2996 8676
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 5852 8732 5916 8736
rect 5852 8676 5856 8732
rect 5856 8676 5912 8732
rect 5912 8676 5916 8732
rect 5852 8672 5916 8676
rect 5932 8732 5996 8736
rect 5932 8676 5936 8732
rect 5936 8676 5992 8732
rect 5992 8676 5996 8732
rect 5932 8672 5996 8676
rect 6012 8732 6076 8736
rect 6012 8676 6016 8732
rect 6016 8676 6072 8732
rect 6072 8676 6076 8732
rect 6012 8672 6076 8676
rect 6092 8732 6156 8736
rect 6092 8676 6096 8732
rect 6096 8676 6152 8732
rect 6152 8676 6156 8732
rect 6092 8672 6156 8676
rect 8852 8732 8916 8736
rect 8852 8676 8856 8732
rect 8856 8676 8912 8732
rect 8912 8676 8916 8732
rect 8852 8672 8916 8676
rect 8932 8732 8996 8736
rect 8932 8676 8936 8732
rect 8936 8676 8992 8732
rect 8992 8676 8996 8732
rect 8932 8672 8996 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 11852 8732 11916 8736
rect 11852 8676 11856 8732
rect 11856 8676 11912 8732
rect 11912 8676 11916 8732
rect 11852 8672 11916 8676
rect 11932 8732 11996 8736
rect 11932 8676 11936 8732
rect 11936 8676 11992 8732
rect 11992 8676 11996 8732
rect 11932 8672 11996 8676
rect 12012 8732 12076 8736
rect 12012 8676 12016 8732
rect 12016 8676 12072 8732
rect 12072 8676 12076 8732
rect 12012 8672 12076 8676
rect 12092 8732 12156 8736
rect 12092 8676 12096 8732
rect 12096 8676 12152 8732
rect 12152 8676 12156 8732
rect 12092 8672 12156 8676
rect 14852 8732 14916 8736
rect 14852 8676 14856 8732
rect 14856 8676 14912 8732
rect 14912 8676 14916 8732
rect 14852 8672 14916 8676
rect 14932 8732 14996 8736
rect 14932 8676 14936 8732
rect 14936 8676 14992 8732
rect 14992 8676 14996 8732
rect 14932 8672 14996 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 17932 8732 17996 8736
rect 17932 8676 17936 8732
rect 17936 8676 17992 8732
rect 17992 8676 17996 8732
rect 17932 8672 17996 8676
rect 18012 8732 18076 8736
rect 18012 8676 18016 8732
rect 18016 8676 18072 8732
rect 18072 8676 18076 8732
rect 18012 8672 18076 8676
rect 18092 8732 18156 8736
rect 18092 8676 18096 8732
rect 18096 8676 18152 8732
rect 18152 8676 18156 8732
rect 18092 8672 18156 8676
rect 20852 8732 20916 8736
rect 20852 8676 20856 8732
rect 20856 8676 20912 8732
rect 20912 8676 20916 8732
rect 20852 8672 20916 8676
rect 20932 8732 20996 8736
rect 20932 8676 20936 8732
rect 20936 8676 20992 8732
rect 20992 8676 20996 8732
rect 20932 8672 20996 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 23852 8732 23916 8736
rect 23852 8676 23856 8732
rect 23856 8676 23912 8732
rect 23912 8676 23916 8732
rect 23852 8672 23916 8676
rect 23932 8732 23996 8736
rect 23932 8676 23936 8732
rect 23936 8676 23992 8732
rect 23992 8676 23996 8732
rect 23932 8672 23996 8676
rect 24012 8732 24076 8736
rect 24012 8676 24016 8732
rect 24016 8676 24072 8732
rect 24072 8676 24076 8732
rect 24012 8672 24076 8676
rect 24092 8732 24156 8736
rect 24092 8676 24096 8732
rect 24096 8676 24152 8732
rect 24152 8676 24156 8732
rect 24092 8672 24156 8676
rect 1352 8188 1416 8192
rect 1352 8132 1356 8188
rect 1356 8132 1412 8188
rect 1412 8132 1416 8188
rect 1352 8128 1416 8132
rect 1432 8188 1496 8192
rect 1432 8132 1436 8188
rect 1436 8132 1492 8188
rect 1492 8132 1496 8188
rect 1432 8128 1496 8132
rect 1512 8188 1576 8192
rect 1512 8132 1516 8188
rect 1516 8132 1572 8188
rect 1572 8132 1576 8188
rect 1512 8128 1576 8132
rect 1592 8188 1656 8192
rect 1592 8132 1596 8188
rect 1596 8132 1652 8188
rect 1652 8132 1656 8188
rect 1592 8128 1656 8132
rect 4352 8188 4416 8192
rect 4352 8132 4356 8188
rect 4356 8132 4412 8188
rect 4412 8132 4416 8188
rect 4352 8128 4416 8132
rect 4432 8188 4496 8192
rect 4432 8132 4436 8188
rect 4436 8132 4492 8188
rect 4492 8132 4496 8188
rect 4432 8128 4496 8132
rect 4512 8188 4576 8192
rect 4512 8132 4516 8188
rect 4516 8132 4572 8188
rect 4572 8132 4576 8188
rect 4512 8128 4576 8132
rect 4592 8188 4656 8192
rect 4592 8132 4596 8188
rect 4596 8132 4652 8188
rect 4652 8132 4656 8188
rect 4592 8128 4656 8132
rect 7352 8188 7416 8192
rect 7352 8132 7356 8188
rect 7356 8132 7412 8188
rect 7412 8132 7416 8188
rect 7352 8128 7416 8132
rect 7432 8188 7496 8192
rect 7432 8132 7436 8188
rect 7436 8132 7492 8188
rect 7492 8132 7496 8188
rect 7432 8128 7496 8132
rect 7512 8188 7576 8192
rect 7512 8132 7516 8188
rect 7516 8132 7572 8188
rect 7572 8132 7576 8188
rect 7512 8128 7576 8132
rect 7592 8188 7656 8192
rect 7592 8132 7596 8188
rect 7596 8132 7652 8188
rect 7652 8132 7656 8188
rect 7592 8128 7656 8132
rect 10352 8188 10416 8192
rect 10352 8132 10356 8188
rect 10356 8132 10412 8188
rect 10412 8132 10416 8188
rect 10352 8128 10416 8132
rect 10432 8188 10496 8192
rect 10432 8132 10436 8188
rect 10436 8132 10492 8188
rect 10492 8132 10496 8188
rect 10432 8128 10496 8132
rect 10512 8188 10576 8192
rect 10512 8132 10516 8188
rect 10516 8132 10572 8188
rect 10572 8132 10576 8188
rect 10512 8128 10576 8132
rect 10592 8188 10656 8192
rect 10592 8132 10596 8188
rect 10596 8132 10652 8188
rect 10652 8132 10656 8188
rect 10592 8128 10656 8132
rect 13352 8188 13416 8192
rect 13352 8132 13356 8188
rect 13356 8132 13412 8188
rect 13412 8132 13416 8188
rect 13352 8128 13416 8132
rect 13432 8188 13496 8192
rect 13432 8132 13436 8188
rect 13436 8132 13492 8188
rect 13492 8132 13496 8188
rect 13432 8128 13496 8132
rect 13512 8188 13576 8192
rect 13512 8132 13516 8188
rect 13516 8132 13572 8188
rect 13572 8132 13576 8188
rect 13512 8128 13576 8132
rect 13592 8188 13656 8192
rect 13592 8132 13596 8188
rect 13596 8132 13652 8188
rect 13652 8132 13656 8188
rect 13592 8128 13656 8132
rect 16352 8188 16416 8192
rect 16352 8132 16356 8188
rect 16356 8132 16412 8188
rect 16412 8132 16416 8188
rect 16352 8128 16416 8132
rect 16432 8188 16496 8192
rect 16432 8132 16436 8188
rect 16436 8132 16492 8188
rect 16492 8132 16496 8188
rect 16432 8128 16496 8132
rect 16512 8188 16576 8192
rect 16512 8132 16516 8188
rect 16516 8132 16572 8188
rect 16572 8132 16576 8188
rect 16512 8128 16576 8132
rect 16592 8188 16656 8192
rect 16592 8132 16596 8188
rect 16596 8132 16652 8188
rect 16652 8132 16656 8188
rect 16592 8128 16656 8132
rect 19352 8188 19416 8192
rect 19352 8132 19356 8188
rect 19356 8132 19412 8188
rect 19412 8132 19416 8188
rect 19352 8128 19416 8132
rect 19432 8188 19496 8192
rect 19432 8132 19436 8188
rect 19436 8132 19492 8188
rect 19492 8132 19496 8188
rect 19432 8128 19496 8132
rect 19512 8188 19576 8192
rect 19512 8132 19516 8188
rect 19516 8132 19572 8188
rect 19572 8132 19576 8188
rect 19512 8128 19576 8132
rect 19592 8188 19656 8192
rect 19592 8132 19596 8188
rect 19596 8132 19652 8188
rect 19652 8132 19656 8188
rect 19592 8128 19656 8132
rect 22352 8188 22416 8192
rect 22352 8132 22356 8188
rect 22356 8132 22412 8188
rect 22412 8132 22416 8188
rect 22352 8128 22416 8132
rect 22432 8188 22496 8192
rect 22432 8132 22436 8188
rect 22436 8132 22492 8188
rect 22492 8132 22496 8188
rect 22432 8128 22496 8132
rect 22512 8188 22576 8192
rect 22512 8132 22516 8188
rect 22516 8132 22572 8188
rect 22572 8132 22576 8188
rect 22512 8128 22576 8132
rect 22592 8188 22656 8192
rect 22592 8132 22596 8188
rect 22596 8132 22652 8188
rect 22652 8132 22656 8188
rect 22592 8128 22656 8132
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 2932 7644 2996 7648
rect 2932 7588 2936 7644
rect 2936 7588 2992 7644
rect 2992 7588 2996 7644
rect 2932 7584 2996 7588
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 5852 7644 5916 7648
rect 5852 7588 5856 7644
rect 5856 7588 5912 7644
rect 5912 7588 5916 7644
rect 5852 7584 5916 7588
rect 5932 7644 5996 7648
rect 5932 7588 5936 7644
rect 5936 7588 5992 7644
rect 5992 7588 5996 7644
rect 5932 7584 5996 7588
rect 6012 7644 6076 7648
rect 6012 7588 6016 7644
rect 6016 7588 6072 7644
rect 6072 7588 6076 7644
rect 6012 7584 6076 7588
rect 6092 7644 6156 7648
rect 6092 7588 6096 7644
rect 6096 7588 6152 7644
rect 6152 7588 6156 7644
rect 6092 7584 6156 7588
rect 8852 7644 8916 7648
rect 8852 7588 8856 7644
rect 8856 7588 8912 7644
rect 8912 7588 8916 7644
rect 8852 7584 8916 7588
rect 8932 7644 8996 7648
rect 8932 7588 8936 7644
rect 8936 7588 8992 7644
rect 8992 7588 8996 7644
rect 8932 7584 8996 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 11852 7644 11916 7648
rect 11852 7588 11856 7644
rect 11856 7588 11912 7644
rect 11912 7588 11916 7644
rect 11852 7584 11916 7588
rect 11932 7644 11996 7648
rect 11932 7588 11936 7644
rect 11936 7588 11992 7644
rect 11992 7588 11996 7644
rect 11932 7584 11996 7588
rect 12012 7644 12076 7648
rect 12012 7588 12016 7644
rect 12016 7588 12072 7644
rect 12072 7588 12076 7644
rect 12012 7584 12076 7588
rect 12092 7644 12156 7648
rect 12092 7588 12096 7644
rect 12096 7588 12152 7644
rect 12152 7588 12156 7644
rect 12092 7584 12156 7588
rect 14852 7644 14916 7648
rect 14852 7588 14856 7644
rect 14856 7588 14912 7644
rect 14912 7588 14916 7644
rect 14852 7584 14916 7588
rect 14932 7644 14996 7648
rect 14932 7588 14936 7644
rect 14936 7588 14992 7644
rect 14992 7588 14996 7644
rect 14932 7584 14996 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 17932 7644 17996 7648
rect 17932 7588 17936 7644
rect 17936 7588 17992 7644
rect 17992 7588 17996 7644
rect 17932 7584 17996 7588
rect 18012 7644 18076 7648
rect 18012 7588 18016 7644
rect 18016 7588 18072 7644
rect 18072 7588 18076 7644
rect 18012 7584 18076 7588
rect 18092 7644 18156 7648
rect 18092 7588 18096 7644
rect 18096 7588 18152 7644
rect 18152 7588 18156 7644
rect 18092 7584 18156 7588
rect 20852 7644 20916 7648
rect 20852 7588 20856 7644
rect 20856 7588 20912 7644
rect 20912 7588 20916 7644
rect 20852 7584 20916 7588
rect 20932 7644 20996 7648
rect 20932 7588 20936 7644
rect 20936 7588 20992 7644
rect 20992 7588 20996 7644
rect 20932 7584 20996 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 23852 7644 23916 7648
rect 23852 7588 23856 7644
rect 23856 7588 23912 7644
rect 23912 7588 23916 7644
rect 23852 7584 23916 7588
rect 23932 7644 23996 7648
rect 23932 7588 23936 7644
rect 23936 7588 23992 7644
rect 23992 7588 23996 7644
rect 23932 7584 23996 7588
rect 24012 7644 24076 7648
rect 24012 7588 24016 7644
rect 24016 7588 24072 7644
rect 24072 7588 24076 7644
rect 24012 7584 24076 7588
rect 24092 7644 24156 7648
rect 24092 7588 24096 7644
rect 24096 7588 24152 7644
rect 24152 7588 24156 7644
rect 24092 7584 24156 7588
rect 1352 7100 1416 7104
rect 1352 7044 1356 7100
rect 1356 7044 1412 7100
rect 1412 7044 1416 7100
rect 1352 7040 1416 7044
rect 1432 7100 1496 7104
rect 1432 7044 1436 7100
rect 1436 7044 1492 7100
rect 1492 7044 1496 7100
rect 1432 7040 1496 7044
rect 1512 7100 1576 7104
rect 1512 7044 1516 7100
rect 1516 7044 1572 7100
rect 1572 7044 1576 7100
rect 1512 7040 1576 7044
rect 1592 7100 1656 7104
rect 1592 7044 1596 7100
rect 1596 7044 1652 7100
rect 1652 7044 1656 7100
rect 1592 7040 1656 7044
rect 4352 7100 4416 7104
rect 4352 7044 4356 7100
rect 4356 7044 4412 7100
rect 4412 7044 4416 7100
rect 4352 7040 4416 7044
rect 4432 7100 4496 7104
rect 4432 7044 4436 7100
rect 4436 7044 4492 7100
rect 4492 7044 4496 7100
rect 4432 7040 4496 7044
rect 4512 7100 4576 7104
rect 4512 7044 4516 7100
rect 4516 7044 4572 7100
rect 4572 7044 4576 7100
rect 4512 7040 4576 7044
rect 4592 7100 4656 7104
rect 4592 7044 4596 7100
rect 4596 7044 4652 7100
rect 4652 7044 4656 7100
rect 4592 7040 4656 7044
rect 7352 7100 7416 7104
rect 7352 7044 7356 7100
rect 7356 7044 7412 7100
rect 7412 7044 7416 7100
rect 7352 7040 7416 7044
rect 7432 7100 7496 7104
rect 7432 7044 7436 7100
rect 7436 7044 7492 7100
rect 7492 7044 7496 7100
rect 7432 7040 7496 7044
rect 7512 7100 7576 7104
rect 7512 7044 7516 7100
rect 7516 7044 7572 7100
rect 7572 7044 7576 7100
rect 7512 7040 7576 7044
rect 7592 7100 7656 7104
rect 7592 7044 7596 7100
rect 7596 7044 7652 7100
rect 7652 7044 7656 7100
rect 7592 7040 7656 7044
rect 10352 7100 10416 7104
rect 10352 7044 10356 7100
rect 10356 7044 10412 7100
rect 10412 7044 10416 7100
rect 10352 7040 10416 7044
rect 10432 7100 10496 7104
rect 10432 7044 10436 7100
rect 10436 7044 10492 7100
rect 10492 7044 10496 7100
rect 10432 7040 10496 7044
rect 10512 7100 10576 7104
rect 10512 7044 10516 7100
rect 10516 7044 10572 7100
rect 10572 7044 10576 7100
rect 10512 7040 10576 7044
rect 10592 7100 10656 7104
rect 10592 7044 10596 7100
rect 10596 7044 10652 7100
rect 10652 7044 10656 7100
rect 10592 7040 10656 7044
rect 13352 7100 13416 7104
rect 13352 7044 13356 7100
rect 13356 7044 13412 7100
rect 13412 7044 13416 7100
rect 13352 7040 13416 7044
rect 13432 7100 13496 7104
rect 13432 7044 13436 7100
rect 13436 7044 13492 7100
rect 13492 7044 13496 7100
rect 13432 7040 13496 7044
rect 13512 7100 13576 7104
rect 13512 7044 13516 7100
rect 13516 7044 13572 7100
rect 13572 7044 13576 7100
rect 13512 7040 13576 7044
rect 13592 7100 13656 7104
rect 13592 7044 13596 7100
rect 13596 7044 13652 7100
rect 13652 7044 13656 7100
rect 13592 7040 13656 7044
rect 16352 7100 16416 7104
rect 16352 7044 16356 7100
rect 16356 7044 16412 7100
rect 16412 7044 16416 7100
rect 16352 7040 16416 7044
rect 16432 7100 16496 7104
rect 16432 7044 16436 7100
rect 16436 7044 16492 7100
rect 16492 7044 16496 7100
rect 16432 7040 16496 7044
rect 16512 7100 16576 7104
rect 16512 7044 16516 7100
rect 16516 7044 16572 7100
rect 16572 7044 16576 7100
rect 16512 7040 16576 7044
rect 16592 7100 16656 7104
rect 16592 7044 16596 7100
rect 16596 7044 16652 7100
rect 16652 7044 16656 7100
rect 16592 7040 16656 7044
rect 19352 7100 19416 7104
rect 19352 7044 19356 7100
rect 19356 7044 19412 7100
rect 19412 7044 19416 7100
rect 19352 7040 19416 7044
rect 19432 7100 19496 7104
rect 19432 7044 19436 7100
rect 19436 7044 19492 7100
rect 19492 7044 19496 7100
rect 19432 7040 19496 7044
rect 19512 7100 19576 7104
rect 19512 7044 19516 7100
rect 19516 7044 19572 7100
rect 19572 7044 19576 7100
rect 19512 7040 19576 7044
rect 19592 7100 19656 7104
rect 19592 7044 19596 7100
rect 19596 7044 19652 7100
rect 19652 7044 19656 7100
rect 19592 7040 19656 7044
rect 22352 7100 22416 7104
rect 22352 7044 22356 7100
rect 22356 7044 22412 7100
rect 22412 7044 22416 7100
rect 22352 7040 22416 7044
rect 22432 7100 22496 7104
rect 22432 7044 22436 7100
rect 22436 7044 22492 7100
rect 22492 7044 22496 7100
rect 22432 7040 22496 7044
rect 22512 7100 22576 7104
rect 22512 7044 22516 7100
rect 22516 7044 22572 7100
rect 22572 7044 22576 7100
rect 22512 7040 22576 7044
rect 22592 7100 22656 7104
rect 22592 7044 22596 7100
rect 22596 7044 22652 7100
rect 22652 7044 22656 7100
rect 22592 7040 22656 7044
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 2932 6556 2996 6560
rect 2932 6500 2936 6556
rect 2936 6500 2992 6556
rect 2992 6500 2996 6556
rect 2932 6496 2996 6500
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 5852 6556 5916 6560
rect 5852 6500 5856 6556
rect 5856 6500 5912 6556
rect 5912 6500 5916 6556
rect 5852 6496 5916 6500
rect 5932 6556 5996 6560
rect 5932 6500 5936 6556
rect 5936 6500 5992 6556
rect 5992 6500 5996 6556
rect 5932 6496 5996 6500
rect 6012 6556 6076 6560
rect 6012 6500 6016 6556
rect 6016 6500 6072 6556
rect 6072 6500 6076 6556
rect 6012 6496 6076 6500
rect 6092 6556 6156 6560
rect 6092 6500 6096 6556
rect 6096 6500 6152 6556
rect 6152 6500 6156 6556
rect 6092 6496 6156 6500
rect 8852 6556 8916 6560
rect 8852 6500 8856 6556
rect 8856 6500 8912 6556
rect 8912 6500 8916 6556
rect 8852 6496 8916 6500
rect 8932 6556 8996 6560
rect 8932 6500 8936 6556
rect 8936 6500 8992 6556
rect 8992 6500 8996 6556
rect 8932 6496 8996 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 11852 6556 11916 6560
rect 11852 6500 11856 6556
rect 11856 6500 11912 6556
rect 11912 6500 11916 6556
rect 11852 6496 11916 6500
rect 11932 6556 11996 6560
rect 11932 6500 11936 6556
rect 11936 6500 11992 6556
rect 11992 6500 11996 6556
rect 11932 6496 11996 6500
rect 12012 6556 12076 6560
rect 12012 6500 12016 6556
rect 12016 6500 12072 6556
rect 12072 6500 12076 6556
rect 12012 6496 12076 6500
rect 12092 6556 12156 6560
rect 12092 6500 12096 6556
rect 12096 6500 12152 6556
rect 12152 6500 12156 6556
rect 12092 6496 12156 6500
rect 14852 6556 14916 6560
rect 14852 6500 14856 6556
rect 14856 6500 14912 6556
rect 14912 6500 14916 6556
rect 14852 6496 14916 6500
rect 14932 6556 14996 6560
rect 14932 6500 14936 6556
rect 14936 6500 14992 6556
rect 14992 6500 14996 6556
rect 14932 6496 14996 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 17932 6556 17996 6560
rect 17932 6500 17936 6556
rect 17936 6500 17992 6556
rect 17992 6500 17996 6556
rect 17932 6496 17996 6500
rect 18012 6556 18076 6560
rect 18012 6500 18016 6556
rect 18016 6500 18072 6556
rect 18072 6500 18076 6556
rect 18012 6496 18076 6500
rect 18092 6556 18156 6560
rect 18092 6500 18096 6556
rect 18096 6500 18152 6556
rect 18152 6500 18156 6556
rect 18092 6496 18156 6500
rect 20852 6556 20916 6560
rect 20852 6500 20856 6556
rect 20856 6500 20912 6556
rect 20912 6500 20916 6556
rect 20852 6496 20916 6500
rect 20932 6556 20996 6560
rect 20932 6500 20936 6556
rect 20936 6500 20992 6556
rect 20992 6500 20996 6556
rect 20932 6496 20996 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 23852 6556 23916 6560
rect 23852 6500 23856 6556
rect 23856 6500 23912 6556
rect 23912 6500 23916 6556
rect 23852 6496 23916 6500
rect 23932 6556 23996 6560
rect 23932 6500 23936 6556
rect 23936 6500 23992 6556
rect 23992 6500 23996 6556
rect 23932 6496 23996 6500
rect 24012 6556 24076 6560
rect 24012 6500 24016 6556
rect 24016 6500 24072 6556
rect 24072 6500 24076 6556
rect 24012 6496 24076 6500
rect 24092 6556 24156 6560
rect 24092 6500 24096 6556
rect 24096 6500 24152 6556
rect 24152 6500 24156 6556
rect 24092 6496 24156 6500
rect 1352 6012 1416 6016
rect 1352 5956 1356 6012
rect 1356 5956 1412 6012
rect 1412 5956 1416 6012
rect 1352 5952 1416 5956
rect 1432 6012 1496 6016
rect 1432 5956 1436 6012
rect 1436 5956 1492 6012
rect 1492 5956 1496 6012
rect 1432 5952 1496 5956
rect 1512 6012 1576 6016
rect 1512 5956 1516 6012
rect 1516 5956 1572 6012
rect 1572 5956 1576 6012
rect 1512 5952 1576 5956
rect 1592 6012 1656 6016
rect 1592 5956 1596 6012
rect 1596 5956 1652 6012
rect 1652 5956 1656 6012
rect 1592 5952 1656 5956
rect 4352 6012 4416 6016
rect 4352 5956 4356 6012
rect 4356 5956 4412 6012
rect 4412 5956 4416 6012
rect 4352 5952 4416 5956
rect 4432 6012 4496 6016
rect 4432 5956 4436 6012
rect 4436 5956 4492 6012
rect 4492 5956 4496 6012
rect 4432 5952 4496 5956
rect 4512 6012 4576 6016
rect 4512 5956 4516 6012
rect 4516 5956 4572 6012
rect 4572 5956 4576 6012
rect 4512 5952 4576 5956
rect 4592 6012 4656 6016
rect 4592 5956 4596 6012
rect 4596 5956 4652 6012
rect 4652 5956 4656 6012
rect 4592 5952 4656 5956
rect 7352 6012 7416 6016
rect 7352 5956 7356 6012
rect 7356 5956 7412 6012
rect 7412 5956 7416 6012
rect 7352 5952 7416 5956
rect 7432 6012 7496 6016
rect 7432 5956 7436 6012
rect 7436 5956 7492 6012
rect 7492 5956 7496 6012
rect 7432 5952 7496 5956
rect 7512 6012 7576 6016
rect 7512 5956 7516 6012
rect 7516 5956 7572 6012
rect 7572 5956 7576 6012
rect 7512 5952 7576 5956
rect 7592 6012 7656 6016
rect 7592 5956 7596 6012
rect 7596 5956 7652 6012
rect 7652 5956 7656 6012
rect 7592 5952 7656 5956
rect 10352 6012 10416 6016
rect 10352 5956 10356 6012
rect 10356 5956 10412 6012
rect 10412 5956 10416 6012
rect 10352 5952 10416 5956
rect 10432 6012 10496 6016
rect 10432 5956 10436 6012
rect 10436 5956 10492 6012
rect 10492 5956 10496 6012
rect 10432 5952 10496 5956
rect 10512 6012 10576 6016
rect 10512 5956 10516 6012
rect 10516 5956 10572 6012
rect 10572 5956 10576 6012
rect 10512 5952 10576 5956
rect 10592 6012 10656 6016
rect 10592 5956 10596 6012
rect 10596 5956 10652 6012
rect 10652 5956 10656 6012
rect 10592 5952 10656 5956
rect 13352 6012 13416 6016
rect 13352 5956 13356 6012
rect 13356 5956 13412 6012
rect 13412 5956 13416 6012
rect 13352 5952 13416 5956
rect 13432 6012 13496 6016
rect 13432 5956 13436 6012
rect 13436 5956 13492 6012
rect 13492 5956 13496 6012
rect 13432 5952 13496 5956
rect 13512 6012 13576 6016
rect 13512 5956 13516 6012
rect 13516 5956 13572 6012
rect 13572 5956 13576 6012
rect 13512 5952 13576 5956
rect 13592 6012 13656 6016
rect 13592 5956 13596 6012
rect 13596 5956 13652 6012
rect 13652 5956 13656 6012
rect 13592 5952 13656 5956
rect 16352 6012 16416 6016
rect 16352 5956 16356 6012
rect 16356 5956 16412 6012
rect 16412 5956 16416 6012
rect 16352 5952 16416 5956
rect 16432 6012 16496 6016
rect 16432 5956 16436 6012
rect 16436 5956 16492 6012
rect 16492 5956 16496 6012
rect 16432 5952 16496 5956
rect 16512 6012 16576 6016
rect 16512 5956 16516 6012
rect 16516 5956 16572 6012
rect 16572 5956 16576 6012
rect 16512 5952 16576 5956
rect 16592 6012 16656 6016
rect 16592 5956 16596 6012
rect 16596 5956 16652 6012
rect 16652 5956 16656 6012
rect 16592 5952 16656 5956
rect 19352 6012 19416 6016
rect 19352 5956 19356 6012
rect 19356 5956 19412 6012
rect 19412 5956 19416 6012
rect 19352 5952 19416 5956
rect 19432 6012 19496 6016
rect 19432 5956 19436 6012
rect 19436 5956 19492 6012
rect 19492 5956 19496 6012
rect 19432 5952 19496 5956
rect 19512 6012 19576 6016
rect 19512 5956 19516 6012
rect 19516 5956 19572 6012
rect 19572 5956 19576 6012
rect 19512 5952 19576 5956
rect 19592 6012 19656 6016
rect 19592 5956 19596 6012
rect 19596 5956 19652 6012
rect 19652 5956 19656 6012
rect 19592 5952 19656 5956
rect 22352 6012 22416 6016
rect 22352 5956 22356 6012
rect 22356 5956 22412 6012
rect 22412 5956 22416 6012
rect 22352 5952 22416 5956
rect 22432 6012 22496 6016
rect 22432 5956 22436 6012
rect 22436 5956 22492 6012
rect 22492 5956 22496 6012
rect 22432 5952 22496 5956
rect 22512 6012 22576 6016
rect 22512 5956 22516 6012
rect 22516 5956 22572 6012
rect 22572 5956 22576 6012
rect 22512 5952 22576 5956
rect 22592 6012 22656 6016
rect 22592 5956 22596 6012
rect 22596 5956 22652 6012
rect 22652 5956 22656 6012
rect 22592 5952 22656 5956
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 2932 5468 2996 5472
rect 2932 5412 2936 5468
rect 2936 5412 2992 5468
rect 2992 5412 2996 5468
rect 2932 5408 2996 5412
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 5852 5468 5916 5472
rect 5852 5412 5856 5468
rect 5856 5412 5912 5468
rect 5912 5412 5916 5468
rect 5852 5408 5916 5412
rect 5932 5468 5996 5472
rect 5932 5412 5936 5468
rect 5936 5412 5992 5468
rect 5992 5412 5996 5468
rect 5932 5408 5996 5412
rect 6012 5468 6076 5472
rect 6012 5412 6016 5468
rect 6016 5412 6072 5468
rect 6072 5412 6076 5468
rect 6012 5408 6076 5412
rect 6092 5468 6156 5472
rect 6092 5412 6096 5468
rect 6096 5412 6152 5468
rect 6152 5412 6156 5468
rect 6092 5408 6156 5412
rect 8852 5468 8916 5472
rect 8852 5412 8856 5468
rect 8856 5412 8912 5468
rect 8912 5412 8916 5468
rect 8852 5408 8916 5412
rect 8932 5468 8996 5472
rect 8932 5412 8936 5468
rect 8936 5412 8992 5468
rect 8992 5412 8996 5468
rect 8932 5408 8996 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 11852 5468 11916 5472
rect 11852 5412 11856 5468
rect 11856 5412 11912 5468
rect 11912 5412 11916 5468
rect 11852 5408 11916 5412
rect 11932 5468 11996 5472
rect 11932 5412 11936 5468
rect 11936 5412 11992 5468
rect 11992 5412 11996 5468
rect 11932 5408 11996 5412
rect 12012 5468 12076 5472
rect 12012 5412 12016 5468
rect 12016 5412 12072 5468
rect 12072 5412 12076 5468
rect 12012 5408 12076 5412
rect 12092 5468 12156 5472
rect 12092 5412 12096 5468
rect 12096 5412 12152 5468
rect 12152 5412 12156 5468
rect 12092 5408 12156 5412
rect 14852 5468 14916 5472
rect 14852 5412 14856 5468
rect 14856 5412 14912 5468
rect 14912 5412 14916 5468
rect 14852 5408 14916 5412
rect 14932 5468 14996 5472
rect 14932 5412 14936 5468
rect 14936 5412 14992 5468
rect 14992 5412 14996 5468
rect 14932 5408 14996 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 17932 5468 17996 5472
rect 17932 5412 17936 5468
rect 17936 5412 17992 5468
rect 17992 5412 17996 5468
rect 17932 5408 17996 5412
rect 18012 5468 18076 5472
rect 18012 5412 18016 5468
rect 18016 5412 18072 5468
rect 18072 5412 18076 5468
rect 18012 5408 18076 5412
rect 18092 5468 18156 5472
rect 18092 5412 18096 5468
rect 18096 5412 18152 5468
rect 18152 5412 18156 5468
rect 18092 5408 18156 5412
rect 20852 5468 20916 5472
rect 20852 5412 20856 5468
rect 20856 5412 20912 5468
rect 20912 5412 20916 5468
rect 20852 5408 20916 5412
rect 20932 5468 20996 5472
rect 20932 5412 20936 5468
rect 20936 5412 20992 5468
rect 20992 5412 20996 5468
rect 20932 5408 20996 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 23852 5468 23916 5472
rect 23852 5412 23856 5468
rect 23856 5412 23912 5468
rect 23912 5412 23916 5468
rect 23852 5408 23916 5412
rect 23932 5468 23996 5472
rect 23932 5412 23936 5468
rect 23936 5412 23992 5468
rect 23992 5412 23996 5468
rect 23932 5408 23996 5412
rect 24012 5468 24076 5472
rect 24012 5412 24016 5468
rect 24016 5412 24072 5468
rect 24072 5412 24076 5468
rect 24012 5408 24076 5412
rect 24092 5468 24156 5472
rect 24092 5412 24096 5468
rect 24096 5412 24152 5468
rect 24152 5412 24156 5468
rect 24092 5408 24156 5412
rect 1352 4924 1416 4928
rect 1352 4868 1356 4924
rect 1356 4868 1412 4924
rect 1412 4868 1416 4924
rect 1352 4864 1416 4868
rect 1432 4924 1496 4928
rect 1432 4868 1436 4924
rect 1436 4868 1492 4924
rect 1492 4868 1496 4924
rect 1432 4864 1496 4868
rect 1512 4924 1576 4928
rect 1512 4868 1516 4924
rect 1516 4868 1572 4924
rect 1572 4868 1576 4924
rect 1512 4864 1576 4868
rect 1592 4924 1656 4928
rect 1592 4868 1596 4924
rect 1596 4868 1652 4924
rect 1652 4868 1656 4924
rect 1592 4864 1656 4868
rect 4352 4924 4416 4928
rect 4352 4868 4356 4924
rect 4356 4868 4412 4924
rect 4412 4868 4416 4924
rect 4352 4864 4416 4868
rect 4432 4924 4496 4928
rect 4432 4868 4436 4924
rect 4436 4868 4492 4924
rect 4492 4868 4496 4924
rect 4432 4864 4496 4868
rect 4512 4924 4576 4928
rect 4512 4868 4516 4924
rect 4516 4868 4572 4924
rect 4572 4868 4576 4924
rect 4512 4864 4576 4868
rect 4592 4924 4656 4928
rect 4592 4868 4596 4924
rect 4596 4868 4652 4924
rect 4652 4868 4656 4924
rect 4592 4864 4656 4868
rect 7352 4924 7416 4928
rect 7352 4868 7356 4924
rect 7356 4868 7412 4924
rect 7412 4868 7416 4924
rect 7352 4864 7416 4868
rect 7432 4924 7496 4928
rect 7432 4868 7436 4924
rect 7436 4868 7492 4924
rect 7492 4868 7496 4924
rect 7432 4864 7496 4868
rect 7512 4924 7576 4928
rect 7512 4868 7516 4924
rect 7516 4868 7572 4924
rect 7572 4868 7576 4924
rect 7512 4864 7576 4868
rect 7592 4924 7656 4928
rect 7592 4868 7596 4924
rect 7596 4868 7652 4924
rect 7652 4868 7656 4924
rect 7592 4864 7656 4868
rect 10352 4924 10416 4928
rect 10352 4868 10356 4924
rect 10356 4868 10412 4924
rect 10412 4868 10416 4924
rect 10352 4864 10416 4868
rect 10432 4924 10496 4928
rect 10432 4868 10436 4924
rect 10436 4868 10492 4924
rect 10492 4868 10496 4924
rect 10432 4864 10496 4868
rect 10512 4924 10576 4928
rect 10512 4868 10516 4924
rect 10516 4868 10572 4924
rect 10572 4868 10576 4924
rect 10512 4864 10576 4868
rect 10592 4924 10656 4928
rect 10592 4868 10596 4924
rect 10596 4868 10652 4924
rect 10652 4868 10656 4924
rect 10592 4864 10656 4868
rect 13352 4924 13416 4928
rect 13352 4868 13356 4924
rect 13356 4868 13412 4924
rect 13412 4868 13416 4924
rect 13352 4864 13416 4868
rect 13432 4924 13496 4928
rect 13432 4868 13436 4924
rect 13436 4868 13492 4924
rect 13492 4868 13496 4924
rect 13432 4864 13496 4868
rect 13512 4924 13576 4928
rect 13512 4868 13516 4924
rect 13516 4868 13572 4924
rect 13572 4868 13576 4924
rect 13512 4864 13576 4868
rect 13592 4924 13656 4928
rect 13592 4868 13596 4924
rect 13596 4868 13652 4924
rect 13652 4868 13656 4924
rect 13592 4864 13656 4868
rect 16352 4924 16416 4928
rect 16352 4868 16356 4924
rect 16356 4868 16412 4924
rect 16412 4868 16416 4924
rect 16352 4864 16416 4868
rect 16432 4924 16496 4928
rect 16432 4868 16436 4924
rect 16436 4868 16492 4924
rect 16492 4868 16496 4924
rect 16432 4864 16496 4868
rect 16512 4924 16576 4928
rect 16512 4868 16516 4924
rect 16516 4868 16572 4924
rect 16572 4868 16576 4924
rect 16512 4864 16576 4868
rect 16592 4924 16656 4928
rect 16592 4868 16596 4924
rect 16596 4868 16652 4924
rect 16652 4868 16656 4924
rect 16592 4864 16656 4868
rect 19352 4924 19416 4928
rect 19352 4868 19356 4924
rect 19356 4868 19412 4924
rect 19412 4868 19416 4924
rect 19352 4864 19416 4868
rect 19432 4924 19496 4928
rect 19432 4868 19436 4924
rect 19436 4868 19492 4924
rect 19492 4868 19496 4924
rect 19432 4864 19496 4868
rect 19512 4924 19576 4928
rect 19512 4868 19516 4924
rect 19516 4868 19572 4924
rect 19572 4868 19576 4924
rect 19512 4864 19576 4868
rect 19592 4924 19656 4928
rect 19592 4868 19596 4924
rect 19596 4868 19652 4924
rect 19652 4868 19656 4924
rect 19592 4864 19656 4868
rect 22352 4924 22416 4928
rect 22352 4868 22356 4924
rect 22356 4868 22412 4924
rect 22412 4868 22416 4924
rect 22352 4864 22416 4868
rect 22432 4924 22496 4928
rect 22432 4868 22436 4924
rect 22436 4868 22492 4924
rect 22492 4868 22496 4924
rect 22432 4864 22496 4868
rect 22512 4924 22576 4928
rect 22512 4868 22516 4924
rect 22516 4868 22572 4924
rect 22572 4868 22576 4924
rect 22512 4864 22576 4868
rect 22592 4924 22656 4928
rect 22592 4868 22596 4924
rect 22596 4868 22652 4924
rect 22652 4868 22656 4924
rect 22592 4864 22656 4868
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 2932 4380 2996 4384
rect 2932 4324 2936 4380
rect 2936 4324 2992 4380
rect 2992 4324 2996 4380
rect 2932 4320 2996 4324
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 5852 4380 5916 4384
rect 5852 4324 5856 4380
rect 5856 4324 5912 4380
rect 5912 4324 5916 4380
rect 5852 4320 5916 4324
rect 5932 4380 5996 4384
rect 5932 4324 5936 4380
rect 5936 4324 5992 4380
rect 5992 4324 5996 4380
rect 5932 4320 5996 4324
rect 6012 4380 6076 4384
rect 6012 4324 6016 4380
rect 6016 4324 6072 4380
rect 6072 4324 6076 4380
rect 6012 4320 6076 4324
rect 6092 4380 6156 4384
rect 6092 4324 6096 4380
rect 6096 4324 6152 4380
rect 6152 4324 6156 4380
rect 6092 4320 6156 4324
rect 8852 4380 8916 4384
rect 8852 4324 8856 4380
rect 8856 4324 8912 4380
rect 8912 4324 8916 4380
rect 8852 4320 8916 4324
rect 8932 4380 8996 4384
rect 8932 4324 8936 4380
rect 8936 4324 8992 4380
rect 8992 4324 8996 4380
rect 8932 4320 8996 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 11852 4380 11916 4384
rect 11852 4324 11856 4380
rect 11856 4324 11912 4380
rect 11912 4324 11916 4380
rect 11852 4320 11916 4324
rect 11932 4380 11996 4384
rect 11932 4324 11936 4380
rect 11936 4324 11992 4380
rect 11992 4324 11996 4380
rect 11932 4320 11996 4324
rect 12012 4380 12076 4384
rect 12012 4324 12016 4380
rect 12016 4324 12072 4380
rect 12072 4324 12076 4380
rect 12012 4320 12076 4324
rect 12092 4380 12156 4384
rect 12092 4324 12096 4380
rect 12096 4324 12152 4380
rect 12152 4324 12156 4380
rect 12092 4320 12156 4324
rect 14852 4380 14916 4384
rect 14852 4324 14856 4380
rect 14856 4324 14912 4380
rect 14912 4324 14916 4380
rect 14852 4320 14916 4324
rect 14932 4380 14996 4384
rect 14932 4324 14936 4380
rect 14936 4324 14992 4380
rect 14992 4324 14996 4380
rect 14932 4320 14996 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 17932 4380 17996 4384
rect 17932 4324 17936 4380
rect 17936 4324 17992 4380
rect 17992 4324 17996 4380
rect 17932 4320 17996 4324
rect 18012 4380 18076 4384
rect 18012 4324 18016 4380
rect 18016 4324 18072 4380
rect 18072 4324 18076 4380
rect 18012 4320 18076 4324
rect 18092 4380 18156 4384
rect 18092 4324 18096 4380
rect 18096 4324 18152 4380
rect 18152 4324 18156 4380
rect 18092 4320 18156 4324
rect 20852 4380 20916 4384
rect 20852 4324 20856 4380
rect 20856 4324 20912 4380
rect 20912 4324 20916 4380
rect 20852 4320 20916 4324
rect 20932 4380 20996 4384
rect 20932 4324 20936 4380
rect 20936 4324 20992 4380
rect 20992 4324 20996 4380
rect 20932 4320 20996 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 23852 4380 23916 4384
rect 23852 4324 23856 4380
rect 23856 4324 23912 4380
rect 23912 4324 23916 4380
rect 23852 4320 23916 4324
rect 23932 4380 23996 4384
rect 23932 4324 23936 4380
rect 23936 4324 23992 4380
rect 23992 4324 23996 4380
rect 23932 4320 23996 4324
rect 24012 4380 24076 4384
rect 24012 4324 24016 4380
rect 24016 4324 24072 4380
rect 24072 4324 24076 4380
rect 24012 4320 24076 4324
rect 24092 4380 24156 4384
rect 24092 4324 24096 4380
rect 24096 4324 24152 4380
rect 24152 4324 24156 4380
rect 24092 4320 24156 4324
rect 1352 3836 1416 3840
rect 1352 3780 1356 3836
rect 1356 3780 1412 3836
rect 1412 3780 1416 3836
rect 1352 3776 1416 3780
rect 1432 3836 1496 3840
rect 1432 3780 1436 3836
rect 1436 3780 1492 3836
rect 1492 3780 1496 3836
rect 1432 3776 1496 3780
rect 1512 3836 1576 3840
rect 1512 3780 1516 3836
rect 1516 3780 1572 3836
rect 1572 3780 1576 3836
rect 1512 3776 1576 3780
rect 1592 3836 1656 3840
rect 1592 3780 1596 3836
rect 1596 3780 1652 3836
rect 1652 3780 1656 3836
rect 1592 3776 1656 3780
rect 4352 3836 4416 3840
rect 4352 3780 4356 3836
rect 4356 3780 4412 3836
rect 4412 3780 4416 3836
rect 4352 3776 4416 3780
rect 4432 3836 4496 3840
rect 4432 3780 4436 3836
rect 4436 3780 4492 3836
rect 4492 3780 4496 3836
rect 4432 3776 4496 3780
rect 4512 3836 4576 3840
rect 4512 3780 4516 3836
rect 4516 3780 4572 3836
rect 4572 3780 4576 3836
rect 4512 3776 4576 3780
rect 4592 3836 4656 3840
rect 4592 3780 4596 3836
rect 4596 3780 4652 3836
rect 4652 3780 4656 3836
rect 4592 3776 4656 3780
rect 7352 3836 7416 3840
rect 7352 3780 7356 3836
rect 7356 3780 7412 3836
rect 7412 3780 7416 3836
rect 7352 3776 7416 3780
rect 7432 3836 7496 3840
rect 7432 3780 7436 3836
rect 7436 3780 7492 3836
rect 7492 3780 7496 3836
rect 7432 3776 7496 3780
rect 7512 3836 7576 3840
rect 7512 3780 7516 3836
rect 7516 3780 7572 3836
rect 7572 3780 7576 3836
rect 7512 3776 7576 3780
rect 7592 3836 7656 3840
rect 7592 3780 7596 3836
rect 7596 3780 7652 3836
rect 7652 3780 7656 3836
rect 7592 3776 7656 3780
rect 10352 3836 10416 3840
rect 10352 3780 10356 3836
rect 10356 3780 10412 3836
rect 10412 3780 10416 3836
rect 10352 3776 10416 3780
rect 10432 3836 10496 3840
rect 10432 3780 10436 3836
rect 10436 3780 10492 3836
rect 10492 3780 10496 3836
rect 10432 3776 10496 3780
rect 10512 3836 10576 3840
rect 10512 3780 10516 3836
rect 10516 3780 10572 3836
rect 10572 3780 10576 3836
rect 10512 3776 10576 3780
rect 10592 3836 10656 3840
rect 10592 3780 10596 3836
rect 10596 3780 10652 3836
rect 10652 3780 10656 3836
rect 10592 3776 10656 3780
rect 13352 3836 13416 3840
rect 13352 3780 13356 3836
rect 13356 3780 13412 3836
rect 13412 3780 13416 3836
rect 13352 3776 13416 3780
rect 13432 3836 13496 3840
rect 13432 3780 13436 3836
rect 13436 3780 13492 3836
rect 13492 3780 13496 3836
rect 13432 3776 13496 3780
rect 13512 3836 13576 3840
rect 13512 3780 13516 3836
rect 13516 3780 13572 3836
rect 13572 3780 13576 3836
rect 13512 3776 13576 3780
rect 13592 3836 13656 3840
rect 13592 3780 13596 3836
rect 13596 3780 13652 3836
rect 13652 3780 13656 3836
rect 13592 3776 13656 3780
rect 16352 3836 16416 3840
rect 16352 3780 16356 3836
rect 16356 3780 16412 3836
rect 16412 3780 16416 3836
rect 16352 3776 16416 3780
rect 16432 3836 16496 3840
rect 16432 3780 16436 3836
rect 16436 3780 16492 3836
rect 16492 3780 16496 3836
rect 16432 3776 16496 3780
rect 16512 3836 16576 3840
rect 16512 3780 16516 3836
rect 16516 3780 16572 3836
rect 16572 3780 16576 3836
rect 16512 3776 16576 3780
rect 16592 3836 16656 3840
rect 16592 3780 16596 3836
rect 16596 3780 16652 3836
rect 16652 3780 16656 3836
rect 16592 3776 16656 3780
rect 19352 3836 19416 3840
rect 19352 3780 19356 3836
rect 19356 3780 19412 3836
rect 19412 3780 19416 3836
rect 19352 3776 19416 3780
rect 19432 3836 19496 3840
rect 19432 3780 19436 3836
rect 19436 3780 19492 3836
rect 19492 3780 19496 3836
rect 19432 3776 19496 3780
rect 19512 3836 19576 3840
rect 19512 3780 19516 3836
rect 19516 3780 19572 3836
rect 19572 3780 19576 3836
rect 19512 3776 19576 3780
rect 19592 3836 19656 3840
rect 19592 3780 19596 3836
rect 19596 3780 19652 3836
rect 19652 3780 19656 3836
rect 19592 3776 19656 3780
rect 22352 3836 22416 3840
rect 22352 3780 22356 3836
rect 22356 3780 22412 3836
rect 22412 3780 22416 3836
rect 22352 3776 22416 3780
rect 22432 3836 22496 3840
rect 22432 3780 22436 3836
rect 22436 3780 22492 3836
rect 22492 3780 22496 3836
rect 22432 3776 22496 3780
rect 22512 3836 22576 3840
rect 22512 3780 22516 3836
rect 22516 3780 22572 3836
rect 22572 3780 22576 3836
rect 22512 3776 22576 3780
rect 22592 3836 22656 3840
rect 22592 3780 22596 3836
rect 22596 3780 22652 3836
rect 22652 3780 22656 3836
rect 22592 3776 22656 3780
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 2932 3292 2996 3296
rect 2932 3236 2936 3292
rect 2936 3236 2992 3292
rect 2992 3236 2996 3292
rect 2932 3232 2996 3236
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 5852 3292 5916 3296
rect 5852 3236 5856 3292
rect 5856 3236 5912 3292
rect 5912 3236 5916 3292
rect 5852 3232 5916 3236
rect 5932 3292 5996 3296
rect 5932 3236 5936 3292
rect 5936 3236 5992 3292
rect 5992 3236 5996 3292
rect 5932 3232 5996 3236
rect 6012 3292 6076 3296
rect 6012 3236 6016 3292
rect 6016 3236 6072 3292
rect 6072 3236 6076 3292
rect 6012 3232 6076 3236
rect 6092 3292 6156 3296
rect 6092 3236 6096 3292
rect 6096 3236 6152 3292
rect 6152 3236 6156 3292
rect 6092 3232 6156 3236
rect 8852 3292 8916 3296
rect 8852 3236 8856 3292
rect 8856 3236 8912 3292
rect 8912 3236 8916 3292
rect 8852 3232 8916 3236
rect 8932 3292 8996 3296
rect 8932 3236 8936 3292
rect 8936 3236 8992 3292
rect 8992 3236 8996 3292
rect 8932 3232 8996 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 11852 3292 11916 3296
rect 11852 3236 11856 3292
rect 11856 3236 11912 3292
rect 11912 3236 11916 3292
rect 11852 3232 11916 3236
rect 11932 3292 11996 3296
rect 11932 3236 11936 3292
rect 11936 3236 11992 3292
rect 11992 3236 11996 3292
rect 11932 3232 11996 3236
rect 12012 3292 12076 3296
rect 12012 3236 12016 3292
rect 12016 3236 12072 3292
rect 12072 3236 12076 3292
rect 12012 3232 12076 3236
rect 12092 3292 12156 3296
rect 12092 3236 12096 3292
rect 12096 3236 12152 3292
rect 12152 3236 12156 3292
rect 12092 3232 12156 3236
rect 14852 3292 14916 3296
rect 14852 3236 14856 3292
rect 14856 3236 14912 3292
rect 14912 3236 14916 3292
rect 14852 3232 14916 3236
rect 14932 3292 14996 3296
rect 14932 3236 14936 3292
rect 14936 3236 14992 3292
rect 14992 3236 14996 3292
rect 14932 3232 14996 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 17932 3292 17996 3296
rect 17932 3236 17936 3292
rect 17936 3236 17992 3292
rect 17992 3236 17996 3292
rect 17932 3232 17996 3236
rect 18012 3292 18076 3296
rect 18012 3236 18016 3292
rect 18016 3236 18072 3292
rect 18072 3236 18076 3292
rect 18012 3232 18076 3236
rect 18092 3292 18156 3296
rect 18092 3236 18096 3292
rect 18096 3236 18152 3292
rect 18152 3236 18156 3292
rect 18092 3232 18156 3236
rect 20852 3292 20916 3296
rect 20852 3236 20856 3292
rect 20856 3236 20912 3292
rect 20912 3236 20916 3292
rect 20852 3232 20916 3236
rect 20932 3292 20996 3296
rect 20932 3236 20936 3292
rect 20936 3236 20992 3292
rect 20992 3236 20996 3292
rect 20932 3232 20996 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 23852 3292 23916 3296
rect 23852 3236 23856 3292
rect 23856 3236 23912 3292
rect 23912 3236 23916 3292
rect 23852 3232 23916 3236
rect 23932 3292 23996 3296
rect 23932 3236 23936 3292
rect 23936 3236 23992 3292
rect 23992 3236 23996 3292
rect 23932 3232 23996 3236
rect 24012 3292 24076 3296
rect 24012 3236 24016 3292
rect 24016 3236 24072 3292
rect 24072 3236 24076 3292
rect 24012 3232 24076 3236
rect 24092 3292 24156 3296
rect 24092 3236 24096 3292
rect 24096 3236 24152 3292
rect 24152 3236 24156 3292
rect 24092 3232 24156 3236
rect 1352 2748 1416 2752
rect 1352 2692 1356 2748
rect 1356 2692 1412 2748
rect 1412 2692 1416 2748
rect 1352 2688 1416 2692
rect 1432 2748 1496 2752
rect 1432 2692 1436 2748
rect 1436 2692 1492 2748
rect 1492 2692 1496 2748
rect 1432 2688 1496 2692
rect 1512 2748 1576 2752
rect 1512 2692 1516 2748
rect 1516 2692 1572 2748
rect 1572 2692 1576 2748
rect 1512 2688 1576 2692
rect 1592 2748 1656 2752
rect 1592 2692 1596 2748
rect 1596 2692 1652 2748
rect 1652 2692 1656 2748
rect 1592 2688 1656 2692
rect 4352 2748 4416 2752
rect 4352 2692 4356 2748
rect 4356 2692 4412 2748
rect 4412 2692 4416 2748
rect 4352 2688 4416 2692
rect 4432 2748 4496 2752
rect 4432 2692 4436 2748
rect 4436 2692 4492 2748
rect 4492 2692 4496 2748
rect 4432 2688 4496 2692
rect 4512 2748 4576 2752
rect 4512 2692 4516 2748
rect 4516 2692 4572 2748
rect 4572 2692 4576 2748
rect 4512 2688 4576 2692
rect 4592 2748 4656 2752
rect 4592 2692 4596 2748
rect 4596 2692 4652 2748
rect 4652 2692 4656 2748
rect 4592 2688 4656 2692
rect 7352 2748 7416 2752
rect 7352 2692 7356 2748
rect 7356 2692 7412 2748
rect 7412 2692 7416 2748
rect 7352 2688 7416 2692
rect 7432 2748 7496 2752
rect 7432 2692 7436 2748
rect 7436 2692 7492 2748
rect 7492 2692 7496 2748
rect 7432 2688 7496 2692
rect 7512 2748 7576 2752
rect 7512 2692 7516 2748
rect 7516 2692 7572 2748
rect 7572 2692 7576 2748
rect 7512 2688 7576 2692
rect 7592 2748 7656 2752
rect 7592 2692 7596 2748
rect 7596 2692 7652 2748
rect 7652 2692 7656 2748
rect 7592 2688 7656 2692
rect 10352 2748 10416 2752
rect 10352 2692 10356 2748
rect 10356 2692 10412 2748
rect 10412 2692 10416 2748
rect 10352 2688 10416 2692
rect 10432 2748 10496 2752
rect 10432 2692 10436 2748
rect 10436 2692 10492 2748
rect 10492 2692 10496 2748
rect 10432 2688 10496 2692
rect 10512 2748 10576 2752
rect 10512 2692 10516 2748
rect 10516 2692 10572 2748
rect 10572 2692 10576 2748
rect 10512 2688 10576 2692
rect 10592 2748 10656 2752
rect 10592 2692 10596 2748
rect 10596 2692 10652 2748
rect 10652 2692 10656 2748
rect 10592 2688 10656 2692
rect 13352 2748 13416 2752
rect 13352 2692 13356 2748
rect 13356 2692 13412 2748
rect 13412 2692 13416 2748
rect 13352 2688 13416 2692
rect 13432 2748 13496 2752
rect 13432 2692 13436 2748
rect 13436 2692 13492 2748
rect 13492 2692 13496 2748
rect 13432 2688 13496 2692
rect 13512 2748 13576 2752
rect 13512 2692 13516 2748
rect 13516 2692 13572 2748
rect 13572 2692 13576 2748
rect 13512 2688 13576 2692
rect 13592 2748 13656 2752
rect 13592 2692 13596 2748
rect 13596 2692 13652 2748
rect 13652 2692 13656 2748
rect 13592 2688 13656 2692
rect 16352 2748 16416 2752
rect 16352 2692 16356 2748
rect 16356 2692 16412 2748
rect 16412 2692 16416 2748
rect 16352 2688 16416 2692
rect 16432 2748 16496 2752
rect 16432 2692 16436 2748
rect 16436 2692 16492 2748
rect 16492 2692 16496 2748
rect 16432 2688 16496 2692
rect 16512 2748 16576 2752
rect 16512 2692 16516 2748
rect 16516 2692 16572 2748
rect 16572 2692 16576 2748
rect 16512 2688 16576 2692
rect 16592 2748 16656 2752
rect 16592 2692 16596 2748
rect 16596 2692 16652 2748
rect 16652 2692 16656 2748
rect 16592 2688 16656 2692
rect 19352 2748 19416 2752
rect 19352 2692 19356 2748
rect 19356 2692 19412 2748
rect 19412 2692 19416 2748
rect 19352 2688 19416 2692
rect 19432 2748 19496 2752
rect 19432 2692 19436 2748
rect 19436 2692 19492 2748
rect 19492 2692 19496 2748
rect 19432 2688 19496 2692
rect 19512 2748 19576 2752
rect 19512 2692 19516 2748
rect 19516 2692 19572 2748
rect 19572 2692 19576 2748
rect 19512 2688 19576 2692
rect 19592 2748 19656 2752
rect 19592 2692 19596 2748
rect 19596 2692 19652 2748
rect 19652 2692 19656 2748
rect 19592 2688 19656 2692
rect 22352 2748 22416 2752
rect 22352 2692 22356 2748
rect 22356 2692 22412 2748
rect 22412 2692 22416 2748
rect 22352 2688 22416 2692
rect 22432 2748 22496 2752
rect 22432 2692 22436 2748
rect 22436 2692 22492 2748
rect 22492 2692 22496 2748
rect 22432 2688 22496 2692
rect 22512 2748 22576 2752
rect 22512 2692 22516 2748
rect 22516 2692 22572 2748
rect 22572 2692 22576 2748
rect 22512 2688 22576 2692
rect 22592 2748 22656 2752
rect 22592 2692 22596 2748
rect 22596 2692 22652 2748
rect 22652 2692 22656 2748
rect 22592 2688 22656 2692
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 2932 2204 2996 2208
rect 2932 2148 2936 2204
rect 2936 2148 2992 2204
rect 2992 2148 2996 2204
rect 2932 2144 2996 2148
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 5852 2204 5916 2208
rect 5852 2148 5856 2204
rect 5856 2148 5912 2204
rect 5912 2148 5916 2204
rect 5852 2144 5916 2148
rect 5932 2204 5996 2208
rect 5932 2148 5936 2204
rect 5936 2148 5992 2204
rect 5992 2148 5996 2204
rect 5932 2144 5996 2148
rect 6012 2204 6076 2208
rect 6012 2148 6016 2204
rect 6016 2148 6072 2204
rect 6072 2148 6076 2204
rect 6012 2144 6076 2148
rect 6092 2204 6156 2208
rect 6092 2148 6096 2204
rect 6096 2148 6152 2204
rect 6152 2148 6156 2204
rect 6092 2144 6156 2148
rect 8852 2204 8916 2208
rect 8852 2148 8856 2204
rect 8856 2148 8912 2204
rect 8912 2148 8916 2204
rect 8852 2144 8916 2148
rect 8932 2204 8996 2208
rect 8932 2148 8936 2204
rect 8936 2148 8992 2204
rect 8992 2148 8996 2204
rect 8932 2144 8996 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 11852 2204 11916 2208
rect 11852 2148 11856 2204
rect 11856 2148 11912 2204
rect 11912 2148 11916 2204
rect 11852 2144 11916 2148
rect 11932 2204 11996 2208
rect 11932 2148 11936 2204
rect 11936 2148 11992 2204
rect 11992 2148 11996 2204
rect 11932 2144 11996 2148
rect 12012 2204 12076 2208
rect 12012 2148 12016 2204
rect 12016 2148 12072 2204
rect 12072 2148 12076 2204
rect 12012 2144 12076 2148
rect 12092 2204 12156 2208
rect 12092 2148 12096 2204
rect 12096 2148 12152 2204
rect 12152 2148 12156 2204
rect 12092 2144 12156 2148
rect 14852 2204 14916 2208
rect 14852 2148 14856 2204
rect 14856 2148 14912 2204
rect 14912 2148 14916 2204
rect 14852 2144 14916 2148
rect 14932 2204 14996 2208
rect 14932 2148 14936 2204
rect 14936 2148 14992 2204
rect 14992 2148 14996 2204
rect 14932 2144 14996 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
rect 17932 2204 17996 2208
rect 17932 2148 17936 2204
rect 17936 2148 17992 2204
rect 17992 2148 17996 2204
rect 17932 2144 17996 2148
rect 18012 2204 18076 2208
rect 18012 2148 18016 2204
rect 18016 2148 18072 2204
rect 18072 2148 18076 2204
rect 18012 2144 18076 2148
rect 18092 2204 18156 2208
rect 18092 2148 18096 2204
rect 18096 2148 18152 2204
rect 18152 2148 18156 2204
rect 18092 2144 18156 2148
rect 20852 2204 20916 2208
rect 20852 2148 20856 2204
rect 20856 2148 20912 2204
rect 20912 2148 20916 2204
rect 20852 2144 20916 2148
rect 20932 2204 20996 2208
rect 20932 2148 20936 2204
rect 20936 2148 20992 2204
rect 20992 2148 20996 2204
rect 20932 2144 20996 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 23852 2204 23916 2208
rect 23852 2148 23856 2204
rect 23856 2148 23912 2204
rect 23912 2148 23916 2204
rect 23852 2144 23916 2148
rect 23932 2204 23996 2208
rect 23932 2148 23936 2204
rect 23936 2148 23992 2204
rect 23992 2148 23996 2204
rect 23932 2144 23996 2148
rect 24012 2204 24076 2208
rect 24012 2148 24016 2204
rect 24016 2148 24072 2204
rect 24072 2148 24076 2204
rect 24012 2144 24076 2148
rect 24092 2204 24156 2208
rect 24092 2148 24096 2204
rect 24096 2148 24152 2204
rect 24152 2148 24156 2204
rect 24092 2144 24156 2148
<< metal4 >>
rect 1344 24512 1664 25072
rect 1344 24448 1352 24512
rect 1416 24448 1432 24512
rect 1496 24448 1512 24512
rect 1576 24448 1592 24512
rect 1656 24448 1664 24512
rect 1344 23424 1664 24448
rect 1344 23360 1352 23424
rect 1416 23360 1432 23424
rect 1496 23360 1512 23424
rect 1576 23360 1592 23424
rect 1656 23360 1664 23424
rect 1344 22336 1664 23360
rect 1344 22272 1352 22336
rect 1416 22272 1432 22336
rect 1496 22272 1512 22336
rect 1576 22272 1592 22336
rect 1656 22272 1664 22336
rect 1344 21248 1664 22272
rect 1344 21184 1352 21248
rect 1416 21184 1432 21248
rect 1496 21184 1512 21248
rect 1576 21184 1592 21248
rect 1656 21184 1664 21248
rect 1344 20160 1664 21184
rect 1344 20096 1352 20160
rect 1416 20096 1432 20160
rect 1496 20096 1512 20160
rect 1576 20096 1592 20160
rect 1656 20096 1664 20160
rect 1344 19072 1664 20096
rect 1344 19008 1352 19072
rect 1416 19008 1432 19072
rect 1496 19008 1512 19072
rect 1576 19008 1592 19072
rect 1656 19008 1664 19072
rect 1344 17984 1664 19008
rect 1344 17920 1352 17984
rect 1416 17920 1432 17984
rect 1496 17920 1512 17984
rect 1576 17920 1592 17984
rect 1656 17920 1664 17984
rect 1344 16896 1664 17920
rect 1344 16832 1352 16896
rect 1416 16832 1432 16896
rect 1496 16832 1512 16896
rect 1576 16832 1592 16896
rect 1656 16832 1664 16896
rect 1344 15808 1664 16832
rect 1344 15744 1352 15808
rect 1416 15744 1432 15808
rect 1496 15744 1512 15808
rect 1576 15744 1592 15808
rect 1656 15744 1664 15808
rect 1344 14720 1664 15744
rect 1344 14656 1352 14720
rect 1416 14656 1432 14720
rect 1496 14656 1512 14720
rect 1576 14656 1592 14720
rect 1656 14656 1664 14720
rect 1344 13632 1664 14656
rect 1344 13568 1352 13632
rect 1416 13568 1432 13632
rect 1496 13568 1512 13632
rect 1576 13568 1592 13632
rect 1656 13568 1664 13632
rect 1344 12544 1664 13568
rect 1344 12480 1352 12544
rect 1416 12480 1432 12544
rect 1496 12480 1512 12544
rect 1576 12480 1592 12544
rect 1656 12480 1664 12544
rect 1344 11456 1664 12480
rect 1344 11392 1352 11456
rect 1416 11392 1432 11456
rect 1496 11392 1512 11456
rect 1576 11392 1592 11456
rect 1656 11392 1664 11456
rect 1344 10368 1664 11392
rect 1344 10304 1352 10368
rect 1416 10304 1432 10368
rect 1496 10304 1512 10368
rect 1576 10304 1592 10368
rect 1656 10304 1664 10368
rect 1344 9280 1664 10304
rect 1344 9216 1352 9280
rect 1416 9216 1432 9280
rect 1496 9216 1512 9280
rect 1576 9216 1592 9280
rect 1656 9216 1664 9280
rect 1344 8192 1664 9216
rect 1344 8128 1352 8192
rect 1416 8128 1432 8192
rect 1496 8128 1512 8192
rect 1576 8128 1592 8192
rect 1656 8128 1664 8192
rect 1344 7104 1664 8128
rect 1344 7040 1352 7104
rect 1416 7040 1432 7104
rect 1496 7040 1512 7104
rect 1576 7040 1592 7104
rect 1656 7040 1664 7104
rect 1344 6016 1664 7040
rect 1344 5952 1352 6016
rect 1416 5952 1432 6016
rect 1496 5952 1512 6016
rect 1576 5952 1592 6016
rect 1656 5952 1664 6016
rect 1344 4928 1664 5952
rect 1344 4864 1352 4928
rect 1416 4864 1432 4928
rect 1496 4864 1512 4928
rect 1576 4864 1592 4928
rect 1656 4864 1664 4928
rect 1344 3840 1664 4864
rect 1344 3776 1352 3840
rect 1416 3776 1432 3840
rect 1496 3776 1512 3840
rect 1576 3776 1592 3840
rect 1656 3776 1664 3840
rect 1344 2752 1664 3776
rect 1344 2688 1352 2752
rect 1416 2688 1432 2752
rect 1496 2688 1512 2752
rect 1576 2688 1592 2752
rect 1656 2688 1664 2752
rect 1344 2128 1664 2688
rect 2844 25056 3164 25072
rect 2844 24992 2852 25056
rect 2916 24992 2932 25056
rect 2996 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3164 25056
rect 2844 23968 3164 24992
rect 2844 23904 2852 23968
rect 2916 23904 2932 23968
rect 2996 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3164 23968
rect 2844 22880 3164 23904
rect 4344 24512 4664 25072
rect 4344 24448 4352 24512
rect 4416 24448 4432 24512
rect 4496 24448 4512 24512
rect 4576 24448 4592 24512
rect 4656 24448 4664 24512
rect 4344 23424 4664 24448
rect 4344 23360 4352 23424
rect 4416 23360 4432 23424
rect 4496 23360 4512 23424
rect 4576 23360 4592 23424
rect 4656 23360 4664 23424
rect 3371 23220 3437 23221
rect 3371 23156 3372 23220
rect 3436 23156 3437 23220
rect 3371 23155 3437 23156
rect 2844 22816 2852 22880
rect 2916 22816 2932 22880
rect 2996 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3164 22880
rect 2844 21792 3164 22816
rect 2844 21728 2852 21792
rect 2916 21728 2932 21792
rect 2996 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3164 21792
rect 2844 20704 3164 21728
rect 2844 20640 2852 20704
rect 2916 20640 2932 20704
rect 2996 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3164 20704
rect 2844 19616 3164 20640
rect 2844 19552 2852 19616
rect 2916 19552 2932 19616
rect 2996 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3164 19616
rect 2844 18528 3164 19552
rect 2844 18464 2852 18528
rect 2916 18464 2932 18528
rect 2996 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3164 18528
rect 2844 17440 3164 18464
rect 2844 17376 2852 17440
rect 2916 17376 2932 17440
rect 2996 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3164 17440
rect 2844 16352 3164 17376
rect 2844 16288 2852 16352
rect 2916 16288 2932 16352
rect 2996 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3164 16352
rect 2844 15264 3164 16288
rect 2844 15200 2852 15264
rect 2916 15200 2932 15264
rect 2996 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3164 15264
rect 2844 14176 3164 15200
rect 2844 14112 2852 14176
rect 2916 14112 2932 14176
rect 2996 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3164 14176
rect 2844 13088 3164 14112
rect 3374 13973 3434 23155
rect 4344 22336 4664 23360
rect 4344 22272 4352 22336
rect 4416 22272 4432 22336
rect 4496 22272 4512 22336
rect 4576 22272 4592 22336
rect 4656 22272 4664 22336
rect 4344 21248 4664 22272
rect 4344 21184 4352 21248
rect 4416 21184 4432 21248
rect 4496 21184 4512 21248
rect 4576 21184 4592 21248
rect 4656 21184 4664 21248
rect 4344 20160 4664 21184
rect 4344 20096 4352 20160
rect 4416 20096 4432 20160
rect 4496 20096 4512 20160
rect 4576 20096 4592 20160
rect 4656 20096 4664 20160
rect 4344 19072 4664 20096
rect 4344 19008 4352 19072
rect 4416 19008 4432 19072
rect 4496 19008 4512 19072
rect 4576 19008 4592 19072
rect 4656 19008 4664 19072
rect 4344 17984 4664 19008
rect 4344 17920 4352 17984
rect 4416 17920 4432 17984
rect 4496 17920 4512 17984
rect 4576 17920 4592 17984
rect 4656 17920 4664 17984
rect 4344 16896 4664 17920
rect 4344 16832 4352 16896
rect 4416 16832 4432 16896
rect 4496 16832 4512 16896
rect 4576 16832 4592 16896
rect 4656 16832 4664 16896
rect 4344 15808 4664 16832
rect 4344 15744 4352 15808
rect 4416 15744 4432 15808
rect 4496 15744 4512 15808
rect 4576 15744 4592 15808
rect 4656 15744 4664 15808
rect 4344 14720 4664 15744
rect 4344 14656 4352 14720
rect 4416 14656 4432 14720
rect 4496 14656 4512 14720
rect 4576 14656 4592 14720
rect 4656 14656 4664 14720
rect 3371 13972 3437 13973
rect 3371 13908 3372 13972
rect 3436 13908 3437 13972
rect 3371 13907 3437 13908
rect 2844 13024 2852 13088
rect 2916 13024 2932 13088
rect 2996 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3164 13088
rect 2844 12000 3164 13024
rect 2844 11936 2852 12000
rect 2916 11936 2932 12000
rect 2996 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3164 12000
rect 2844 10912 3164 11936
rect 2844 10848 2852 10912
rect 2916 10848 2932 10912
rect 2996 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3164 10912
rect 2844 9824 3164 10848
rect 2844 9760 2852 9824
rect 2916 9760 2932 9824
rect 2996 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3164 9824
rect 2844 8736 3164 9760
rect 2844 8672 2852 8736
rect 2916 8672 2932 8736
rect 2996 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3164 8736
rect 2844 7648 3164 8672
rect 2844 7584 2852 7648
rect 2916 7584 2932 7648
rect 2996 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3164 7648
rect 2844 6560 3164 7584
rect 2844 6496 2852 6560
rect 2916 6496 2932 6560
rect 2996 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3164 6560
rect 2844 5472 3164 6496
rect 2844 5408 2852 5472
rect 2916 5408 2932 5472
rect 2996 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3164 5472
rect 2844 4384 3164 5408
rect 2844 4320 2852 4384
rect 2916 4320 2932 4384
rect 2996 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3164 4384
rect 2844 3296 3164 4320
rect 2844 3232 2852 3296
rect 2916 3232 2932 3296
rect 2996 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3164 3296
rect 2844 2208 3164 3232
rect 2844 2144 2852 2208
rect 2916 2144 2932 2208
rect 2996 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3164 2208
rect 2844 2128 3164 2144
rect 4344 13632 4664 14656
rect 4344 13568 4352 13632
rect 4416 13568 4432 13632
rect 4496 13568 4512 13632
rect 4576 13568 4592 13632
rect 4656 13568 4664 13632
rect 4344 12544 4664 13568
rect 4344 12480 4352 12544
rect 4416 12480 4432 12544
rect 4496 12480 4512 12544
rect 4576 12480 4592 12544
rect 4656 12480 4664 12544
rect 4344 11456 4664 12480
rect 4344 11392 4352 11456
rect 4416 11392 4432 11456
rect 4496 11392 4512 11456
rect 4576 11392 4592 11456
rect 4656 11392 4664 11456
rect 4344 10368 4664 11392
rect 4344 10304 4352 10368
rect 4416 10304 4432 10368
rect 4496 10304 4512 10368
rect 4576 10304 4592 10368
rect 4656 10304 4664 10368
rect 4344 9280 4664 10304
rect 4344 9216 4352 9280
rect 4416 9216 4432 9280
rect 4496 9216 4512 9280
rect 4576 9216 4592 9280
rect 4656 9216 4664 9280
rect 4344 8192 4664 9216
rect 4344 8128 4352 8192
rect 4416 8128 4432 8192
rect 4496 8128 4512 8192
rect 4576 8128 4592 8192
rect 4656 8128 4664 8192
rect 4344 7104 4664 8128
rect 4344 7040 4352 7104
rect 4416 7040 4432 7104
rect 4496 7040 4512 7104
rect 4576 7040 4592 7104
rect 4656 7040 4664 7104
rect 4344 6016 4664 7040
rect 4344 5952 4352 6016
rect 4416 5952 4432 6016
rect 4496 5952 4512 6016
rect 4576 5952 4592 6016
rect 4656 5952 4664 6016
rect 4344 4928 4664 5952
rect 4344 4864 4352 4928
rect 4416 4864 4432 4928
rect 4496 4864 4512 4928
rect 4576 4864 4592 4928
rect 4656 4864 4664 4928
rect 4344 3840 4664 4864
rect 4344 3776 4352 3840
rect 4416 3776 4432 3840
rect 4496 3776 4512 3840
rect 4576 3776 4592 3840
rect 4656 3776 4664 3840
rect 4344 2752 4664 3776
rect 4344 2688 4352 2752
rect 4416 2688 4432 2752
rect 4496 2688 4512 2752
rect 4576 2688 4592 2752
rect 4656 2688 4664 2752
rect 4344 2128 4664 2688
rect 5844 25056 6164 25072
rect 5844 24992 5852 25056
rect 5916 24992 5932 25056
rect 5996 24992 6012 25056
rect 6076 24992 6092 25056
rect 6156 24992 6164 25056
rect 5844 23968 6164 24992
rect 5844 23904 5852 23968
rect 5916 23904 5932 23968
rect 5996 23904 6012 23968
rect 6076 23904 6092 23968
rect 6156 23904 6164 23968
rect 5844 22880 6164 23904
rect 5844 22816 5852 22880
rect 5916 22816 5932 22880
rect 5996 22816 6012 22880
rect 6076 22816 6092 22880
rect 6156 22816 6164 22880
rect 5844 21792 6164 22816
rect 5844 21728 5852 21792
rect 5916 21728 5932 21792
rect 5996 21728 6012 21792
rect 6076 21728 6092 21792
rect 6156 21728 6164 21792
rect 5844 20704 6164 21728
rect 5844 20640 5852 20704
rect 5916 20640 5932 20704
rect 5996 20640 6012 20704
rect 6076 20640 6092 20704
rect 6156 20640 6164 20704
rect 5844 19616 6164 20640
rect 5844 19552 5852 19616
rect 5916 19552 5932 19616
rect 5996 19552 6012 19616
rect 6076 19552 6092 19616
rect 6156 19552 6164 19616
rect 5844 18528 6164 19552
rect 5844 18464 5852 18528
rect 5916 18464 5932 18528
rect 5996 18464 6012 18528
rect 6076 18464 6092 18528
rect 6156 18464 6164 18528
rect 5844 17440 6164 18464
rect 5844 17376 5852 17440
rect 5916 17376 5932 17440
rect 5996 17376 6012 17440
rect 6076 17376 6092 17440
rect 6156 17376 6164 17440
rect 5844 16352 6164 17376
rect 5844 16288 5852 16352
rect 5916 16288 5932 16352
rect 5996 16288 6012 16352
rect 6076 16288 6092 16352
rect 6156 16288 6164 16352
rect 5844 15264 6164 16288
rect 5844 15200 5852 15264
rect 5916 15200 5932 15264
rect 5996 15200 6012 15264
rect 6076 15200 6092 15264
rect 6156 15200 6164 15264
rect 5844 14176 6164 15200
rect 5844 14112 5852 14176
rect 5916 14112 5932 14176
rect 5996 14112 6012 14176
rect 6076 14112 6092 14176
rect 6156 14112 6164 14176
rect 5844 13088 6164 14112
rect 5844 13024 5852 13088
rect 5916 13024 5932 13088
rect 5996 13024 6012 13088
rect 6076 13024 6092 13088
rect 6156 13024 6164 13088
rect 5844 12000 6164 13024
rect 5844 11936 5852 12000
rect 5916 11936 5932 12000
rect 5996 11936 6012 12000
rect 6076 11936 6092 12000
rect 6156 11936 6164 12000
rect 5844 10912 6164 11936
rect 5844 10848 5852 10912
rect 5916 10848 5932 10912
rect 5996 10848 6012 10912
rect 6076 10848 6092 10912
rect 6156 10848 6164 10912
rect 5844 9824 6164 10848
rect 5844 9760 5852 9824
rect 5916 9760 5932 9824
rect 5996 9760 6012 9824
rect 6076 9760 6092 9824
rect 6156 9760 6164 9824
rect 5844 8736 6164 9760
rect 5844 8672 5852 8736
rect 5916 8672 5932 8736
rect 5996 8672 6012 8736
rect 6076 8672 6092 8736
rect 6156 8672 6164 8736
rect 5844 7648 6164 8672
rect 5844 7584 5852 7648
rect 5916 7584 5932 7648
rect 5996 7584 6012 7648
rect 6076 7584 6092 7648
rect 6156 7584 6164 7648
rect 5844 6560 6164 7584
rect 5844 6496 5852 6560
rect 5916 6496 5932 6560
rect 5996 6496 6012 6560
rect 6076 6496 6092 6560
rect 6156 6496 6164 6560
rect 5844 5472 6164 6496
rect 5844 5408 5852 5472
rect 5916 5408 5932 5472
rect 5996 5408 6012 5472
rect 6076 5408 6092 5472
rect 6156 5408 6164 5472
rect 5844 4384 6164 5408
rect 5844 4320 5852 4384
rect 5916 4320 5932 4384
rect 5996 4320 6012 4384
rect 6076 4320 6092 4384
rect 6156 4320 6164 4384
rect 5844 3296 6164 4320
rect 5844 3232 5852 3296
rect 5916 3232 5932 3296
rect 5996 3232 6012 3296
rect 6076 3232 6092 3296
rect 6156 3232 6164 3296
rect 5844 2208 6164 3232
rect 5844 2144 5852 2208
rect 5916 2144 5932 2208
rect 5996 2144 6012 2208
rect 6076 2144 6092 2208
rect 6156 2144 6164 2208
rect 5844 2128 6164 2144
rect 7344 24512 7664 25072
rect 7344 24448 7352 24512
rect 7416 24448 7432 24512
rect 7496 24448 7512 24512
rect 7576 24448 7592 24512
rect 7656 24448 7664 24512
rect 7344 23424 7664 24448
rect 7344 23360 7352 23424
rect 7416 23360 7432 23424
rect 7496 23360 7512 23424
rect 7576 23360 7592 23424
rect 7656 23360 7664 23424
rect 7344 22336 7664 23360
rect 7344 22272 7352 22336
rect 7416 22272 7432 22336
rect 7496 22272 7512 22336
rect 7576 22272 7592 22336
rect 7656 22272 7664 22336
rect 7344 21248 7664 22272
rect 7344 21184 7352 21248
rect 7416 21184 7432 21248
rect 7496 21184 7512 21248
rect 7576 21184 7592 21248
rect 7656 21184 7664 21248
rect 7344 20160 7664 21184
rect 7344 20096 7352 20160
rect 7416 20096 7432 20160
rect 7496 20096 7512 20160
rect 7576 20096 7592 20160
rect 7656 20096 7664 20160
rect 7344 19072 7664 20096
rect 7344 19008 7352 19072
rect 7416 19008 7432 19072
rect 7496 19008 7512 19072
rect 7576 19008 7592 19072
rect 7656 19008 7664 19072
rect 7344 17984 7664 19008
rect 7344 17920 7352 17984
rect 7416 17920 7432 17984
rect 7496 17920 7512 17984
rect 7576 17920 7592 17984
rect 7656 17920 7664 17984
rect 7344 16896 7664 17920
rect 7344 16832 7352 16896
rect 7416 16832 7432 16896
rect 7496 16832 7512 16896
rect 7576 16832 7592 16896
rect 7656 16832 7664 16896
rect 7344 15808 7664 16832
rect 7344 15744 7352 15808
rect 7416 15744 7432 15808
rect 7496 15744 7512 15808
rect 7576 15744 7592 15808
rect 7656 15744 7664 15808
rect 7344 14720 7664 15744
rect 7344 14656 7352 14720
rect 7416 14656 7432 14720
rect 7496 14656 7512 14720
rect 7576 14656 7592 14720
rect 7656 14656 7664 14720
rect 7344 13632 7664 14656
rect 7344 13568 7352 13632
rect 7416 13568 7432 13632
rect 7496 13568 7512 13632
rect 7576 13568 7592 13632
rect 7656 13568 7664 13632
rect 7344 12544 7664 13568
rect 7344 12480 7352 12544
rect 7416 12480 7432 12544
rect 7496 12480 7512 12544
rect 7576 12480 7592 12544
rect 7656 12480 7664 12544
rect 7344 11456 7664 12480
rect 7344 11392 7352 11456
rect 7416 11392 7432 11456
rect 7496 11392 7512 11456
rect 7576 11392 7592 11456
rect 7656 11392 7664 11456
rect 7344 10368 7664 11392
rect 7344 10304 7352 10368
rect 7416 10304 7432 10368
rect 7496 10304 7512 10368
rect 7576 10304 7592 10368
rect 7656 10304 7664 10368
rect 7344 9280 7664 10304
rect 7344 9216 7352 9280
rect 7416 9216 7432 9280
rect 7496 9216 7512 9280
rect 7576 9216 7592 9280
rect 7656 9216 7664 9280
rect 7344 8192 7664 9216
rect 7344 8128 7352 8192
rect 7416 8128 7432 8192
rect 7496 8128 7512 8192
rect 7576 8128 7592 8192
rect 7656 8128 7664 8192
rect 7344 7104 7664 8128
rect 7344 7040 7352 7104
rect 7416 7040 7432 7104
rect 7496 7040 7512 7104
rect 7576 7040 7592 7104
rect 7656 7040 7664 7104
rect 7344 6016 7664 7040
rect 7344 5952 7352 6016
rect 7416 5952 7432 6016
rect 7496 5952 7512 6016
rect 7576 5952 7592 6016
rect 7656 5952 7664 6016
rect 7344 4928 7664 5952
rect 7344 4864 7352 4928
rect 7416 4864 7432 4928
rect 7496 4864 7512 4928
rect 7576 4864 7592 4928
rect 7656 4864 7664 4928
rect 7344 3840 7664 4864
rect 7344 3776 7352 3840
rect 7416 3776 7432 3840
rect 7496 3776 7512 3840
rect 7576 3776 7592 3840
rect 7656 3776 7664 3840
rect 7344 2752 7664 3776
rect 7344 2688 7352 2752
rect 7416 2688 7432 2752
rect 7496 2688 7512 2752
rect 7576 2688 7592 2752
rect 7656 2688 7664 2752
rect 7344 2128 7664 2688
rect 8844 25056 9164 25072
rect 8844 24992 8852 25056
rect 8916 24992 8932 25056
rect 8996 24992 9012 25056
rect 9076 24992 9092 25056
rect 9156 24992 9164 25056
rect 8844 23968 9164 24992
rect 8844 23904 8852 23968
rect 8916 23904 8932 23968
rect 8996 23904 9012 23968
rect 9076 23904 9092 23968
rect 9156 23904 9164 23968
rect 8844 22880 9164 23904
rect 8844 22816 8852 22880
rect 8916 22816 8932 22880
rect 8996 22816 9012 22880
rect 9076 22816 9092 22880
rect 9156 22816 9164 22880
rect 8844 21792 9164 22816
rect 8844 21728 8852 21792
rect 8916 21728 8932 21792
rect 8996 21728 9012 21792
rect 9076 21728 9092 21792
rect 9156 21728 9164 21792
rect 8844 20704 9164 21728
rect 8844 20640 8852 20704
rect 8916 20640 8932 20704
rect 8996 20640 9012 20704
rect 9076 20640 9092 20704
rect 9156 20640 9164 20704
rect 8844 19616 9164 20640
rect 8844 19552 8852 19616
rect 8916 19552 8932 19616
rect 8996 19552 9012 19616
rect 9076 19552 9092 19616
rect 9156 19552 9164 19616
rect 8844 18528 9164 19552
rect 8844 18464 8852 18528
rect 8916 18464 8932 18528
rect 8996 18464 9012 18528
rect 9076 18464 9092 18528
rect 9156 18464 9164 18528
rect 8844 17440 9164 18464
rect 8844 17376 8852 17440
rect 8916 17376 8932 17440
rect 8996 17376 9012 17440
rect 9076 17376 9092 17440
rect 9156 17376 9164 17440
rect 8844 16352 9164 17376
rect 8844 16288 8852 16352
rect 8916 16288 8932 16352
rect 8996 16288 9012 16352
rect 9076 16288 9092 16352
rect 9156 16288 9164 16352
rect 8844 15264 9164 16288
rect 8844 15200 8852 15264
rect 8916 15200 8932 15264
rect 8996 15200 9012 15264
rect 9076 15200 9092 15264
rect 9156 15200 9164 15264
rect 8844 14176 9164 15200
rect 8844 14112 8852 14176
rect 8916 14112 8932 14176
rect 8996 14112 9012 14176
rect 9076 14112 9092 14176
rect 9156 14112 9164 14176
rect 8844 13088 9164 14112
rect 8844 13024 8852 13088
rect 8916 13024 8932 13088
rect 8996 13024 9012 13088
rect 9076 13024 9092 13088
rect 9156 13024 9164 13088
rect 8844 12000 9164 13024
rect 8844 11936 8852 12000
rect 8916 11936 8932 12000
rect 8996 11936 9012 12000
rect 9076 11936 9092 12000
rect 9156 11936 9164 12000
rect 8844 10912 9164 11936
rect 8844 10848 8852 10912
rect 8916 10848 8932 10912
rect 8996 10848 9012 10912
rect 9076 10848 9092 10912
rect 9156 10848 9164 10912
rect 8844 9824 9164 10848
rect 8844 9760 8852 9824
rect 8916 9760 8932 9824
rect 8996 9760 9012 9824
rect 9076 9760 9092 9824
rect 9156 9760 9164 9824
rect 8844 8736 9164 9760
rect 8844 8672 8852 8736
rect 8916 8672 8932 8736
rect 8996 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9164 8736
rect 8844 7648 9164 8672
rect 8844 7584 8852 7648
rect 8916 7584 8932 7648
rect 8996 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9164 7648
rect 8844 6560 9164 7584
rect 8844 6496 8852 6560
rect 8916 6496 8932 6560
rect 8996 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9164 6560
rect 8844 5472 9164 6496
rect 8844 5408 8852 5472
rect 8916 5408 8932 5472
rect 8996 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9164 5472
rect 8844 4384 9164 5408
rect 8844 4320 8852 4384
rect 8916 4320 8932 4384
rect 8996 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9164 4384
rect 8844 3296 9164 4320
rect 8844 3232 8852 3296
rect 8916 3232 8932 3296
rect 8996 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9164 3296
rect 8844 2208 9164 3232
rect 8844 2144 8852 2208
rect 8916 2144 8932 2208
rect 8996 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9164 2208
rect 8844 2128 9164 2144
rect 10344 24512 10664 25072
rect 10344 24448 10352 24512
rect 10416 24448 10432 24512
rect 10496 24448 10512 24512
rect 10576 24448 10592 24512
rect 10656 24448 10664 24512
rect 10344 23424 10664 24448
rect 10344 23360 10352 23424
rect 10416 23360 10432 23424
rect 10496 23360 10512 23424
rect 10576 23360 10592 23424
rect 10656 23360 10664 23424
rect 10344 22336 10664 23360
rect 10344 22272 10352 22336
rect 10416 22272 10432 22336
rect 10496 22272 10512 22336
rect 10576 22272 10592 22336
rect 10656 22272 10664 22336
rect 10344 21248 10664 22272
rect 10344 21184 10352 21248
rect 10416 21184 10432 21248
rect 10496 21184 10512 21248
rect 10576 21184 10592 21248
rect 10656 21184 10664 21248
rect 10344 20160 10664 21184
rect 10344 20096 10352 20160
rect 10416 20096 10432 20160
rect 10496 20096 10512 20160
rect 10576 20096 10592 20160
rect 10656 20096 10664 20160
rect 10344 19072 10664 20096
rect 10344 19008 10352 19072
rect 10416 19008 10432 19072
rect 10496 19008 10512 19072
rect 10576 19008 10592 19072
rect 10656 19008 10664 19072
rect 10344 17984 10664 19008
rect 10344 17920 10352 17984
rect 10416 17920 10432 17984
rect 10496 17920 10512 17984
rect 10576 17920 10592 17984
rect 10656 17920 10664 17984
rect 10344 16896 10664 17920
rect 10344 16832 10352 16896
rect 10416 16832 10432 16896
rect 10496 16832 10512 16896
rect 10576 16832 10592 16896
rect 10656 16832 10664 16896
rect 10344 15808 10664 16832
rect 10344 15744 10352 15808
rect 10416 15744 10432 15808
rect 10496 15744 10512 15808
rect 10576 15744 10592 15808
rect 10656 15744 10664 15808
rect 10344 14720 10664 15744
rect 10344 14656 10352 14720
rect 10416 14656 10432 14720
rect 10496 14656 10512 14720
rect 10576 14656 10592 14720
rect 10656 14656 10664 14720
rect 10344 13632 10664 14656
rect 10344 13568 10352 13632
rect 10416 13568 10432 13632
rect 10496 13568 10512 13632
rect 10576 13568 10592 13632
rect 10656 13568 10664 13632
rect 10344 12544 10664 13568
rect 10344 12480 10352 12544
rect 10416 12480 10432 12544
rect 10496 12480 10512 12544
rect 10576 12480 10592 12544
rect 10656 12480 10664 12544
rect 10344 11456 10664 12480
rect 10344 11392 10352 11456
rect 10416 11392 10432 11456
rect 10496 11392 10512 11456
rect 10576 11392 10592 11456
rect 10656 11392 10664 11456
rect 10344 10368 10664 11392
rect 10344 10304 10352 10368
rect 10416 10304 10432 10368
rect 10496 10304 10512 10368
rect 10576 10304 10592 10368
rect 10656 10304 10664 10368
rect 10344 9280 10664 10304
rect 10344 9216 10352 9280
rect 10416 9216 10432 9280
rect 10496 9216 10512 9280
rect 10576 9216 10592 9280
rect 10656 9216 10664 9280
rect 10344 8192 10664 9216
rect 10344 8128 10352 8192
rect 10416 8128 10432 8192
rect 10496 8128 10512 8192
rect 10576 8128 10592 8192
rect 10656 8128 10664 8192
rect 10344 7104 10664 8128
rect 10344 7040 10352 7104
rect 10416 7040 10432 7104
rect 10496 7040 10512 7104
rect 10576 7040 10592 7104
rect 10656 7040 10664 7104
rect 10344 6016 10664 7040
rect 10344 5952 10352 6016
rect 10416 5952 10432 6016
rect 10496 5952 10512 6016
rect 10576 5952 10592 6016
rect 10656 5952 10664 6016
rect 10344 4928 10664 5952
rect 10344 4864 10352 4928
rect 10416 4864 10432 4928
rect 10496 4864 10512 4928
rect 10576 4864 10592 4928
rect 10656 4864 10664 4928
rect 10344 3840 10664 4864
rect 10344 3776 10352 3840
rect 10416 3776 10432 3840
rect 10496 3776 10512 3840
rect 10576 3776 10592 3840
rect 10656 3776 10664 3840
rect 10344 2752 10664 3776
rect 10344 2688 10352 2752
rect 10416 2688 10432 2752
rect 10496 2688 10512 2752
rect 10576 2688 10592 2752
rect 10656 2688 10664 2752
rect 10344 2128 10664 2688
rect 11844 25056 12164 25072
rect 11844 24992 11852 25056
rect 11916 24992 11932 25056
rect 11996 24992 12012 25056
rect 12076 24992 12092 25056
rect 12156 24992 12164 25056
rect 11844 23968 12164 24992
rect 11844 23904 11852 23968
rect 11916 23904 11932 23968
rect 11996 23904 12012 23968
rect 12076 23904 12092 23968
rect 12156 23904 12164 23968
rect 11844 22880 12164 23904
rect 11844 22816 11852 22880
rect 11916 22816 11932 22880
rect 11996 22816 12012 22880
rect 12076 22816 12092 22880
rect 12156 22816 12164 22880
rect 11844 21792 12164 22816
rect 11844 21728 11852 21792
rect 11916 21728 11932 21792
rect 11996 21728 12012 21792
rect 12076 21728 12092 21792
rect 12156 21728 12164 21792
rect 11844 20704 12164 21728
rect 11844 20640 11852 20704
rect 11916 20640 11932 20704
rect 11996 20640 12012 20704
rect 12076 20640 12092 20704
rect 12156 20640 12164 20704
rect 11844 19616 12164 20640
rect 11844 19552 11852 19616
rect 11916 19552 11932 19616
rect 11996 19552 12012 19616
rect 12076 19552 12092 19616
rect 12156 19552 12164 19616
rect 11844 18528 12164 19552
rect 11844 18464 11852 18528
rect 11916 18464 11932 18528
rect 11996 18464 12012 18528
rect 12076 18464 12092 18528
rect 12156 18464 12164 18528
rect 11844 17440 12164 18464
rect 13344 24512 13664 25072
rect 13344 24448 13352 24512
rect 13416 24448 13432 24512
rect 13496 24448 13512 24512
rect 13576 24448 13592 24512
rect 13656 24448 13664 24512
rect 13344 23424 13664 24448
rect 13344 23360 13352 23424
rect 13416 23360 13432 23424
rect 13496 23360 13512 23424
rect 13576 23360 13592 23424
rect 13656 23360 13664 23424
rect 13344 22336 13664 23360
rect 13344 22272 13352 22336
rect 13416 22272 13432 22336
rect 13496 22272 13512 22336
rect 13576 22272 13592 22336
rect 13656 22272 13664 22336
rect 13344 21248 13664 22272
rect 13344 21184 13352 21248
rect 13416 21184 13432 21248
rect 13496 21184 13512 21248
rect 13576 21184 13592 21248
rect 13656 21184 13664 21248
rect 13344 20160 13664 21184
rect 13344 20096 13352 20160
rect 13416 20096 13432 20160
rect 13496 20096 13512 20160
rect 13576 20096 13592 20160
rect 13656 20096 13664 20160
rect 13344 19072 13664 20096
rect 13344 19008 13352 19072
rect 13416 19008 13432 19072
rect 13496 19008 13512 19072
rect 13576 19008 13592 19072
rect 13656 19008 13664 19072
rect 13123 18324 13189 18325
rect 13123 18260 13124 18324
rect 13188 18260 13189 18324
rect 13123 18259 13189 18260
rect 11844 17376 11852 17440
rect 11916 17376 11932 17440
rect 11996 17376 12012 17440
rect 12076 17376 12092 17440
rect 12156 17376 12164 17440
rect 11844 16352 12164 17376
rect 11844 16288 11852 16352
rect 11916 16288 11932 16352
rect 11996 16288 12012 16352
rect 12076 16288 12092 16352
rect 12156 16288 12164 16352
rect 11844 15264 12164 16288
rect 11844 15200 11852 15264
rect 11916 15200 11932 15264
rect 11996 15200 12012 15264
rect 12076 15200 12092 15264
rect 12156 15200 12164 15264
rect 11844 14176 12164 15200
rect 11844 14112 11852 14176
rect 11916 14112 11932 14176
rect 11996 14112 12012 14176
rect 12076 14112 12092 14176
rect 12156 14112 12164 14176
rect 11844 13088 12164 14112
rect 13126 13973 13186 18259
rect 13344 17984 13664 19008
rect 13344 17920 13352 17984
rect 13416 17920 13432 17984
rect 13496 17920 13512 17984
rect 13576 17920 13592 17984
rect 13656 17920 13664 17984
rect 13344 16896 13664 17920
rect 13344 16832 13352 16896
rect 13416 16832 13432 16896
rect 13496 16832 13512 16896
rect 13576 16832 13592 16896
rect 13656 16832 13664 16896
rect 13344 15808 13664 16832
rect 13344 15744 13352 15808
rect 13416 15744 13432 15808
rect 13496 15744 13512 15808
rect 13576 15744 13592 15808
rect 13656 15744 13664 15808
rect 13344 14720 13664 15744
rect 13344 14656 13352 14720
rect 13416 14656 13432 14720
rect 13496 14656 13512 14720
rect 13576 14656 13592 14720
rect 13656 14656 13664 14720
rect 13123 13972 13189 13973
rect 13123 13908 13124 13972
rect 13188 13908 13189 13972
rect 13123 13907 13189 13908
rect 11844 13024 11852 13088
rect 11916 13024 11932 13088
rect 11996 13024 12012 13088
rect 12076 13024 12092 13088
rect 12156 13024 12164 13088
rect 11844 12000 12164 13024
rect 11844 11936 11852 12000
rect 11916 11936 11932 12000
rect 11996 11936 12012 12000
rect 12076 11936 12092 12000
rect 12156 11936 12164 12000
rect 11844 10912 12164 11936
rect 13126 11117 13186 13907
rect 13344 13632 13664 14656
rect 13344 13568 13352 13632
rect 13416 13568 13432 13632
rect 13496 13568 13512 13632
rect 13576 13568 13592 13632
rect 13656 13568 13664 13632
rect 13344 12544 13664 13568
rect 13344 12480 13352 12544
rect 13416 12480 13432 12544
rect 13496 12480 13512 12544
rect 13576 12480 13592 12544
rect 13656 12480 13664 12544
rect 13344 11456 13664 12480
rect 13344 11392 13352 11456
rect 13416 11392 13432 11456
rect 13496 11392 13512 11456
rect 13576 11392 13592 11456
rect 13656 11392 13664 11456
rect 13123 11116 13189 11117
rect 13123 11052 13124 11116
rect 13188 11052 13189 11116
rect 13123 11051 13189 11052
rect 11844 10848 11852 10912
rect 11916 10848 11932 10912
rect 11996 10848 12012 10912
rect 12076 10848 12092 10912
rect 12156 10848 12164 10912
rect 11844 9824 12164 10848
rect 11844 9760 11852 9824
rect 11916 9760 11932 9824
rect 11996 9760 12012 9824
rect 12076 9760 12092 9824
rect 12156 9760 12164 9824
rect 11844 8736 12164 9760
rect 11844 8672 11852 8736
rect 11916 8672 11932 8736
rect 11996 8672 12012 8736
rect 12076 8672 12092 8736
rect 12156 8672 12164 8736
rect 11844 7648 12164 8672
rect 11844 7584 11852 7648
rect 11916 7584 11932 7648
rect 11996 7584 12012 7648
rect 12076 7584 12092 7648
rect 12156 7584 12164 7648
rect 11844 6560 12164 7584
rect 11844 6496 11852 6560
rect 11916 6496 11932 6560
rect 11996 6496 12012 6560
rect 12076 6496 12092 6560
rect 12156 6496 12164 6560
rect 11844 5472 12164 6496
rect 11844 5408 11852 5472
rect 11916 5408 11932 5472
rect 11996 5408 12012 5472
rect 12076 5408 12092 5472
rect 12156 5408 12164 5472
rect 11844 4384 12164 5408
rect 11844 4320 11852 4384
rect 11916 4320 11932 4384
rect 11996 4320 12012 4384
rect 12076 4320 12092 4384
rect 12156 4320 12164 4384
rect 11844 3296 12164 4320
rect 11844 3232 11852 3296
rect 11916 3232 11932 3296
rect 11996 3232 12012 3296
rect 12076 3232 12092 3296
rect 12156 3232 12164 3296
rect 11844 2208 12164 3232
rect 11844 2144 11852 2208
rect 11916 2144 11932 2208
rect 11996 2144 12012 2208
rect 12076 2144 12092 2208
rect 12156 2144 12164 2208
rect 11844 2128 12164 2144
rect 13344 10368 13664 11392
rect 13344 10304 13352 10368
rect 13416 10304 13432 10368
rect 13496 10304 13512 10368
rect 13576 10304 13592 10368
rect 13656 10304 13664 10368
rect 13344 9280 13664 10304
rect 13344 9216 13352 9280
rect 13416 9216 13432 9280
rect 13496 9216 13512 9280
rect 13576 9216 13592 9280
rect 13656 9216 13664 9280
rect 13344 8192 13664 9216
rect 13344 8128 13352 8192
rect 13416 8128 13432 8192
rect 13496 8128 13512 8192
rect 13576 8128 13592 8192
rect 13656 8128 13664 8192
rect 13344 7104 13664 8128
rect 13344 7040 13352 7104
rect 13416 7040 13432 7104
rect 13496 7040 13512 7104
rect 13576 7040 13592 7104
rect 13656 7040 13664 7104
rect 13344 6016 13664 7040
rect 13344 5952 13352 6016
rect 13416 5952 13432 6016
rect 13496 5952 13512 6016
rect 13576 5952 13592 6016
rect 13656 5952 13664 6016
rect 13344 4928 13664 5952
rect 13344 4864 13352 4928
rect 13416 4864 13432 4928
rect 13496 4864 13512 4928
rect 13576 4864 13592 4928
rect 13656 4864 13664 4928
rect 13344 3840 13664 4864
rect 13344 3776 13352 3840
rect 13416 3776 13432 3840
rect 13496 3776 13512 3840
rect 13576 3776 13592 3840
rect 13656 3776 13664 3840
rect 13344 2752 13664 3776
rect 13344 2688 13352 2752
rect 13416 2688 13432 2752
rect 13496 2688 13512 2752
rect 13576 2688 13592 2752
rect 13656 2688 13664 2752
rect 13344 2128 13664 2688
rect 14844 25056 15164 25072
rect 14844 24992 14852 25056
rect 14916 24992 14932 25056
rect 14996 24992 15012 25056
rect 15076 24992 15092 25056
rect 15156 24992 15164 25056
rect 14844 23968 15164 24992
rect 14844 23904 14852 23968
rect 14916 23904 14932 23968
rect 14996 23904 15012 23968
rect 15076 23904 15092 23968
rect 15156 23904 15164 23968
rect 14844 22880 15164 23904
rect 14844 22816 14852 22880
rect 14916 22816 14932 22880
rect 14996 22816 15012 22880
rect 15076 22816 15092 22880
rect 15156 22816 15164 22880
rect 14844 21792 15164 22816
rect 14844 21728 14852 21792
rect 14916 21728 14932 21792
rect 14996 21728 15012 21792
rect 15076 21728 15092 21792
rect 15156 21728 15164 21792
rect 14844 20704 15164 21728
rect 14844 20640 14852 20704
rect 14916 20640 14932 20704
rect 14996 20640 15012 20704
rect 15076 20640 15092 20704
rect 15156 20640 15164 20704
rect 14844 19616 15164 20640
rect 14844 19552 14852 19616
rect 14916 19552 14932 19616
rect 14996 19552 15012 19616
rect 15076 19552 15092 19616
rect 15156 19552 15164 19616
rect 14844 18528 15164 19552
rect 14844 18464 14852 18528
rect 14916 18464 14932 18528
rect 14996 18464 15012 18528
rect 15076 18464 15092 18528
rect 15156 18464 15164 18528
rect 14844 17440 15164 18464
rect 14844 17376 14852 17440
rect 14916 17376 14932 17440
rect 14996 17376 15012 17440
rect 15076 17376 15092 17440
rect 15156 17376 15164 17440
rect 14844 16352 15164 17376
rect 14844 16288 14852 16352
rect 14916 16288 14932 16352
rect 14996 16288 15012 16352
rect 15076 16288 15092 16352
rect 15156 16288 15164 16352
rect 14844 15264 15164 16288
rect 14844 15200 14852 15264
rect 14916 15200 14932 15264
rect 14996 15200 15012 15264
rect 15076 15200 15092 15264
rect 15156 15200 15164 15264
rect 14844 14176 15164 15200
rect 14844 14112 14852 14176
rect 14916 14112 14932 14176
rect 14996 14112 15012 14176
rect 15076 14112 15092 14176
rect 15156 14112 15164 14176
rect 14844 13088 15164 14112
rect 14844 13024 14852 13088
rect 14916 13024 14932 13088
rect 14996 13024 15012 13088
rect 15076 13024 15092 13088
rect 15156 13024 15164 13088
rect 14844 12000 15164 13024
rect 14844 11936 14852 12000
rect 14916 11936 14932 12000
rect 14996 11936 15012 12000
rect 15076 11936 15092 12000
rect 15156 11936 15164 12000
rect 14844 10912 15164 11936
rect 14844 10848 14852 10912
rect 14916 10848 14932 10912
rect 14996 10848 15012 10912
rect 15076 10848 15092 10912
rect 15156 10848 15164 10912
rect 14844 9824 15164 10848
rect 14844 9760 14852 9824
rect 14916 9760 14932 9824
rect 14996 9760 15012 9824
rect 15076 9760 15092 9824
rect 15156 9760 15164 9824
rect 14844 8736 15164 9760
rect 14844 8672 14852 8736
rect 14916 8672 14932 8736
rect 14996 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15164 8736
rect 14844 7648 15164 8672
rect 14844 7584 14852 7648
rect 14916 7584 14932 7648
rect 14996 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15164 7648
rect 14844 6560 15164 7584
rect 14844 6496 14852 6560
rect 14916 6496 14932 6560
rect 14996 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15164 6560
rect 14844 5472 15164 6496
rect 14844 5408 14852 5472
rect 14916 5408 14932 5472
rect 14996 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15164 5472
rect 14844 4384 15164 5408
rect 14844 4320 14852 4384
rect 14916 4320 14932 4384
rect 14996 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15164 4384
rect 14844 3296 15164 4320
rect 14844 3232 14852 3296
rect 14916 3232 14932 3296
rect 14996 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15164 3296
rect 14844 2208 15164 3232
rect 14844 2144 14852 2208
rect 14916 2144 14932 2208
rect 14996 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15164 2208
rect 14844 2128 15164 2144
rect 16344 24512 16664 25072
rect 16344 24448 16352 24512
rect 16416 24448 16432 24512
rect 16496 24448 16512 24512
rect 16576 24448 16592 24512
rect 16656 24448 16664 24512
rect 16344 23424 16664 24448
rect 16344 23360 16352 23424
rect 16416 23360 16432 23424
rect 16496 23360 16512 23424
rect 16576 23360 16592 23424
rect 16656 23360 16664 23424
rect 16344 22336 16664 23360
rect 16344 22272 16352 22336
rect 16416 22272 16432 22336
rect 16496 22272 16512 22336
rect 16576 22272 16592 22336
rect 16656 22272 16664 22336
rect 16344 21248 16664 22272
rect 16344 21184 16352 21248
rect 16416 21184 16432 21248
rect 16496 21184 16512 21248
rect 16576 21184 16592 21248
rect 16656 21184 16664 21248
rect 16344 20160 16664 21184
rect 16344 20096 16352 20160
rect 16416 20096 16432 20160
rect 16496 20096 16512 20160
rect 16576 20096 16592 20160
rect 16656 20096 16664 20160
rect 16344 19072 16664 20096
rect 16344 19008 16352 19072
rect 16416 19008 16432 19072
rect 16496 19008 16512 19072
rect 16576 19008 16592 19072
rect 16656 19008 16664 19072
rect 16344 17984 16664 19008
rect 16344 17920 16352 17984
rect 16416 17920 16432 17984
rect 16496 17920 16512 17984
rect 16576 17920 16592 17984
rect 16656 17920 16664 17984
rect 16344 16896 16664 17920
rect 16344 16832 16352 16896
rect 16416 16832 16432 16896
rect 16496 16832 16512 16896
rect 16576 16832 16592 16896
rect 16656 16832 16664 16896
rect 16344 15808 16664 16832
rect 16344 15744 16352 15808
rect 16416 15744 16432 15808
rect 16496 15744 16512 15808
rect 16576 15744 16592 15808
rect 16656 15744 16664 15808
rect 16344 14720 16664 15744
rect 16344 14656 16352 14720
rect 16416 14656 16432 14720
rect 16496 14656 16512 14720
rect 16576 14656 16592 14720
rect 16656 14656 16664 14720
rect 16344 13632 16664 14656
rect 16344 13568 16352 13632
rect 16416 13568 16432 13632
rect 16496 13568 16512 13632
rect 16576 13568 16592 13632
rect 16656 13568 16664 13632
rect 16344 12544 16664 13568
rect 16344 12480 16352 12544
rect 16416 12480 16432 12544
rect 16496 12480 16512 12544
rect 16576 12480 16592 12544
rect 16656 12480 16664 12544
rect 16344 11456 16664 12480
rect 16344 11392 16352 11456
rect 16416 11392 16432 11456
rect 16496 11392 16512 11456
rect 16576 11392 16592 11456
rect 16656 11392 16664 11456
rect 16344 10368 16664 11392
rect 16344 10304 16352 10368
rect 16416 10304 16432 10368
rect 16496 10304 16512 10368
rect 16576 10304 16592 10368
rect 16656 10304 16664 10368
rect 16344 9280 16664 10304
rect 16344 9216 16352 9280
rect 16416 9216 16432 9280
rect 16496 9216 16512 9280
rect 16576 9216 16592 9280
rect 16656 9216 16664 9280
rect 16344 8192 16664 9216
rect 16344 8128 16352 8192
rect 16416 8128 16432 8192
rect 16496 8128 16512 8192
rect 16576 8128 16592 8192
rect 16656 8128 16664 8192
rect 16344 7104 16664 8128
rect 16344 7040 16352 7104
rect 16416 7040 16432 7104
rect 16496 7040 16512 7104
rect 16576 7040 16592 7104
rect 16656 7040 16664 7104
rect 16344 6016 16664 7040
rect 16344 5952 16352 6016
rect 16416 5952 16432 6016
rect 16496 5952 16512 6016
rect 16576 5952 16592 6016
rect 16656 5952 16664 6016
rect 16344 4928 16664 5952
rect 16344 4864 16352 4928
rect 16416 4864 16432 4928
rect 16496 4864 16512 4928
rect 16576 4864 16592 4928
rect 16656 4864 16664 4928
rect 16344 3840 16664 4864
rect 16344 3776 16352 3840
rect 16416 3776 16432 3840
rect 16496 3776 16512 3840
rect 16576 3776 16592 3840
rect 16656 3776 16664 3840
rect 16344 2752 16664 3776
rect 16344 2688 16352 2752
rect 16416 2688 16432 2752
rect 16496 2688 16512 2752
rect 16576 2688 16592 2752
rect 16656 2688 16664 2752
rect 16344 2128 16664 2688
rect 17844 25056 18164 25072
rect 17844 24992 17852 25056
rect 17916 24992 17932 25056
rect 17996 24992 18012 25056
rect 18076 24992 18092 25056
rect 18156 24992 18164 25056
rect 17844 23968 18164 24992
rect 17844 23904 17852 23968
rect 17916 23904 17932 23968
rect 17996 23904 18012 23968
rect 18076 23904 18092 23968
rect 18156 23904 18164 23968
rect 17844 22880 18164 23904
rect 17844 22816 17852 22880
rect 17916 22816 17932 22880
rect 17996 22816 18012 22880
rect 18076 22816 18092 22880
rect 18156 22816 18164 22880
rect 17844 21792 18164 22816
rect 17844 21728 17852 21792
rect 17916 21728 17932 21792
rect 17996 21728 18012 21792
rect 18076 21728 18092 21792
rect 18156 21728 18164 21792
rect 17844 20704 18164 21728
rect 17844 20640 17852 20704
rect 17916 20640 17932 20704
rect 17996 20640 18012 20704
rect 18076 20640 18092 20704
rect 18156 20640 18164 20704
rect 17844 19616 18164 20640
rect 17844 19552 17852 19616
rect 17916 19552 17932 19616
rect 17996 19552 18012 19616
rect 18076 19552 18092 19616
rect 18156 19552 18164 19616
rect 17844 18528 18164 19552
rect 17844 18464 17852 18528
rect 17916 18464 17932 18528
rect 17996 18464 18012 18528
rect 18076 18464 18092 18528
rect 18156 18464 18164 18528
rect 17844 17440 18164 18464
rect 17844 17376 17852 17440
rect 17916 17376 17932 17440
rect 17996 17376 18012 17440
rect 18076 17376 18092 17440
rect 18156 17376 18164 17440
rect 17844 16352 18164 17376
rect 17844 16288 17852 16352
rect 17916 16288 17932 16352
rect 17996 16288 18012 16352
rect 18076 16288 18092 16352
rect 18156 16288 18164 16352
rect 17844 15264 18164 16288
rect 17844 15200 17852 15264
rect 17916 15200 17932 15264
rect 17996 15200 18012 15264
rect 18076 15200 18092 15264
rect 18156 15200 18164 15264
rect 17844 14176 18164 15200
rect 17844 14112 17852 14176
rect 17916 14112 17932 14176
rect 17996 14112 18012 14176
rect 18076 14112 18092 14176
rect 18156 14112 18164 14176
rect 17844 13088 18164 14112
rect 17844 13024 17852 13088
rect 17916 13024 17932 13088
rect 17996 13024 18012 13088
rect 18076 13024 18092 13088
rect 18156 13024 18164 13088
rect 17844 12000 18164 13024
rect 17844 11936 17852 12000
rect 17916 11936 17932 12000
rect 17996 11936 18012 12000
rect 18076 11936 18092 12000
rect 18156 11936 18164 12000
rect 17844 10912 18164 11936
rect 17844 10848 17852 10912
rect 17916 10848 17932 10912
rect 17996 10848 18012 10912
rect 18076 10848 18092 10912
rect 18156 10848 18164 10912
rect 17844 9824 18164 10848
rect 17844 9760 17852 9824
rect 17916 9760 17932 9824
rect 17996 9760 18012 9824
rect 18076 9760 18092 9824
rect 18156 9760 18164 9824
rect 17844 8736 18164 9760
rect 17844 8672 17852 8736
rect 17916 8672 17932 8736
rect 17996 8672 18012 8736
rect 18076 8672 18092 8736
rect 18156 8672 18164 8736
rect 17844 7648 18164 8672
rect 17844 7584 17852 7648
rect 17916 7584 17932 7648
rect 17996 7584 18012 7648
rect 18076 7584 18092 7648
rect 18156 7584 18164 7648
rect 17844 6560 18164 7584
rect 17844 6496 17852 6560
rect 17916 6496 17932 6560
rect 17996 6496 18012 6560
rect 18076 6496 18092 6560
rect 18156 6496 18164 6560
rect 17844 5472 18164 6496
rect 17844 5408 17852 5472
rect 17916 5408 17932 5472
rect 17996 5408 18012 5472
rect 18076 5408 18092 5472
rect 18156 5408 18164 5472
rect 17844 4384 18164 5408
rect 17844 4320 17852 4384
rect 17916 4320 17932 4384
rect 17996 4320 18012 4384
rect 18076 4320 18092 4384
rect 18156 4320 18164 4384
rect 17844 3296 18164 4320
rect 17844 3232 17852 3296
rect 17916 3232 17932 3296
rect 17996 3232 18012 3296
rect 18076 3232 18092 3296
rect 18156 3232 18164 3296
rect 17844 2208 18164 3232
rect 17844 2144 17852 2208
rect 17916 2144 17932 2208
rect 17996 2144 18012 2208
rect 18076 2144 18092 2208
rect 18156 2144 18164 2208
rect 17844 2128 18164 2144
rect 19344 24512 19664 25072
rect 19344 24448 19352 24512
rect 19416 24448 19432 24512
rect 19496 24448 19512 24512
rect 19576 24448 19592 24512
rect 19656 24448 19664 24512
rect 19344 23424 19664 24448
rect 19344 23360 19352 23424
rect 19416 23360 19432 23424
rect 19496 23360 19512 23424
rect 19576 23360 19592 23424
rect 19656 23360 19664 23424
rect 19344 22336 19664 23360
rect 19344 22272 19352 22336
rect 19416 22272 19432 22336
rect 19496 22272 19512 22336
rect 19576 22272 19592 22336
rect 19656 22272 19664 22336
rect 19344 21248 19664 22272
rect 19344 21184 19352 21248
rect 19416 21184 19432 21248
rect 19496 21184 19512 21248
rect 19576 21184 19592 21248
rect 19656 21184 19664 21248
rect 19344 20160 19664 21184
rect 19344 20096 19352 20160
rect 19416 20096 19432 20160
rect 19496 20096 19512 20160
rect 19576 20096 19592 20160
rect 19656 20096 19664 20160
rect 19344 19072 19664 20096
rect 19344 19008 19352 19072
rect 19416 19008 19432 19072
rect 19496 19008 19512 19072
rect 19576 19008 19592 19072
rect 19656 19008 19664 19072
rect 19344 17984 19664 19008
rect 19344 17920 19352 17984
rect 19416 17920 19432 17984
rect 19496 17920 19512 17984
rect 19576 17920 19592 17984
rect 19656 17920 19664 17984
rect 19344 16896 19664 17920
rect 19344 16832 19352 16896
rect 19416 16832 19432 16896
rect 19496 16832 19512 16896
rect 19576 16832 19592 16896
rect 19656 16832 19664 16896
rect 19344 15808 19664 16832
rect 19344 15744 19352 15808
rect 19416 15744 19432 15808
rect 19496 15744 19512 15808
rect 19576 15744 19592 15808
rect 19656 15744 19664 15808
rect 19344 14720 19664 15744
rect 19344 14656 19352 14720
rect 19416 14656 19432 14720
rect 19496 14656 19512 14720
rect 19576 14656 19592 14720
rect 19656 14656 19664 14720
rect 19344 13632 19664 14656
rect 19344 13568 19352 13632
rect 19416 13568 19432 13632
rect 19496 13568 19512 13632
rect 19576 13568 19592 13632
rect 19656 13568 19664 13632
rect 19344 12544 19664 13568
rect 19344 12480 19352 12544
rect 19416 12480 19432 12544
rect 19496 12480 19512 12544
rect 19576 12480 19592 12544
rect 19656 12480 19664 12544
rect 19344 11456 19664 12480
rect 19344 11392 19352 11456
rect 19416 11392 19432 11456
rect 19496 11392 19512 11456
rect 19576 11392 19592 11456
rect 19656 11392 19664 11456
rect 19344 10368 19664 11392
rect 19344 10304 19352 10368
rect 19416 10304 19432 10368
rect 19496 10304 19512 10368
rect 19576 10304 19592 10368
rect 19656 10304 19664 10368
rect 19344 9280 19664 10304
rect 19344 9216 19352 9280
rect 19416 9216 19432 9280
rect 19496 9216 19512 9280
rect 19576 9216 19592 9280
rect 19656 9216 19664 9280
rect 19344 8192 19664 9216
rect 19344 8128 19352 8192
rect 19416 8128 19432 8192
rect 19496 8128 19512 8192
rect 19576 8128 19592 8192
rect 19656 8128 19664 8192
rect 19344 7104 19664 8128
rect 19344 7040 19352 7104
rect 19416 7040 19432 7104
rect 19496 7040 19512 7104
rect 19576 7040 19592 7104
rect 19656 7040 19664 7104
rect 19344 6016 19664 7040
rect 19344 5952 19352 6016
rect 19416 5952 19432 6016
rect 19496 5952 19512 6016
rect 19576 5952 19592 6016
rect 19656 5952 19664 6016
rect 19344 4928 19664 5952
rect 19344 4864 19352 4928
rect 19416 4864 19432 4928
rect 19496 4864 19512 4928
rect 19576 4864 19592 4928
rect 19656 4864 19664 4928
rect 19344 3840 19664 4864
rect 19344 3776 19352 3840
rect 19416 3776 19432 3840
rect 19496 3776 19512 3840
rect 19576 3776 19592 3840
rect 19656 3776 19664 3840
rect 19344 2752 19664 3776
rect 19344 2688 19352 2752
rect 19416 2688 19432 2752
rect 19496 2688 19512 2752
rect 19576 2688 19592 2752
rect 19656 2688 19664 2752
rect 19344 2128 19664 2688
rect 20844 25056 21164 25072
rect 20844 24992 20852 25056
rect 20916 24992 20932 25056
rect 20996 24992 21012 25056
rect 21076 24992 21092 25056
rect 21156 24992 21164 25056
rect 20844 23968 21164 24992
rect 20844 23904 20852 23968
rect 20916 23904 20932 23968
rect 20996 23904 21012 23968
rect 21076 23904 21092 23968
rect 21156 23904 21164 23968
rect 20844 22880 21164 23904
rect 20844 22816 20852 22880
rect 20916 22816 20932 22880
rect 20996 22816 21012 22880
rect 21076 22816 21092 22880
rect 21156 22816 21164 22880
rect 20844 21792 21164 22816
rect 20844 21728 20852 21792
rect 20916 21728 20932 21792
rect 20996 21728 21012 21792
rect 21076 21728 21092 21792
rect 21156 21728 21164 21792
rect 20844 20704 21164 21728
rect 20844 20640 20852 20704
rect 20916 20640 20932 20704
rect 20996 20640 21012 20704
rect 21076 20640 21092 20704
rect 21156 20640 21164 20704
rect 20844 19616 21164 20640
rect 20844 19552 20852 19616
rect 20916 19552 20932 19616
rect 20996 19552 21012 19616
rect 21076 19552 21092 19616
rect 21156 19552 21164 19616
rect 20844 18528 21164 19552
rect 20844 18464 20852 18528
rect 20916 18464 20932 18528
rect 20996 18464 21012 18528
rect 21076 18464 21092 18528
rect 21156 18464 21164 18528
rect 20844 17440 21164 18464
rect 22344 24512 22664 25072
rect 22344 24448 22352 24512
rect 22416 24448 22432 24512
rect 22496 24448 22512 24512
rect 22576 24448 22592 24512
rect 22656 24448 22664 24512
rect 22344 23424 22664 24448
rect 22344 23360 22352 23424
rect 22416 23360 22432 23424
rect 22496 23360 22512 23424
rect 22576 23360 22592 23424
rect 22656 23360 22664 23424
rect 22344 22336 22664 23360
rect 22344 22272 22352 22336
rect 22416 22272 22432 22336
rect 22496 22272 22512 22336
rect 22576 22272 22592 22336
rect 22656 22272 22664 22336
rect 22344 21248 22664 22272
rect 22344 21184 22352 21248
rect 22416 21184 22432 21248
rect 22496 21184 22512 21248
rect 22576 21184 22592 21248
rect 22656 21184 22664 21248
rect 22344 20160 22664 21184
rect 22344 20096 22352 20160
rect 22416 20096 22432 20160
rect 22496 20096 22512 20160
rect 22576 20096 22592 20160
rect 22656 20096 22664 20160
rect 22344 19072 22664 20096
rect 22344 19008 22352 19072
rect 22416 19008 22432 19072
rect 22496 19008 22512 19072
rect 22576 19008 22592 19072
rect 22656 19008 22664 19072
rect 22139 18188 22205 18189
rect 22139 18124 22140 18188
rect 22204 18124 22205 18188
rect 22139 18123 22205 18124
rect 20844 17376 20852 17440
rect 20916 17376 20932 17440
rect 20996 17376 21012 17440
rect 21076 17376 21092 17440
rect 21156 17376 21164 17440
rect 20844 16352 21164 17376
rect 20844 16288 20852 16352
rect 20916 16288 20932 16352
rect 20996 16288 21012 16352
rect 21076 16288 21092 16352
rect 21156 16288 21164 16352
rect 20844 15264 21164 16288
rect 20844 15200 20852 15264
rect 20916 15200 20932 15264
rect 20996 15200 21012 15264
rect 21076 15200 21092 15264
rect 21156 15200 21164 15264
rect 20844 14176 21164 15200
rect 20844 14112 20852 14176
rect 20916 14112 20932 14176
rect 20996 14112 21012 14176
rect 21076 14112 21092 14176
rect 21156 14112 21164 14176
rect 20844 13088 21164 14112
rect 22142 13701 22202 18123
rect 22344 17984 22664 19008
rect 22344 17920 22352 17984
rect 22416 17920 22432 17984
rect 22496 17920 22512 17984
rect 22576 17920 22592 17984
rect 22656 17920 22664 17984
rect 22344 16896 22664 17920
rect 22344 16832 22352 16896
rect 22416 16832 22432 16896
rect 22496 16832 22512 16896
rect 22576 16832 22592 16896
rect 22656 16832 22664 16896
rect 22344 15808 22664 16832
rect 22344 15744 22352 15808
rect 22416 15744 22432 15808
rect 22496 15744 22512 15808
rect 22576 15744 22592 15808
rect 22656 15744 22664 15808
rect 22344 14720 22664 15744
rect 22344 14656 22352 14720
rect 22416 14656 22432 14720
rect 22496 14656 22512 14720
rect 22576 14656 22592 14720
rect 22656 14656 22664 14720
rect 22139 13700 22205 13701
rect 22139 13636 22140 13700
rect 22204 13636 22205 13700
rect 22139 13635 22205 13636
rect 20844 13024 20852 13088
rect 20916 13024 20932 13088
rect 20996 13024 21012 13088
rect 21076 13024 21092 13088
rect 21156 13024 21164 13088
rect 20844 12000 21164 13024
rect 20844 11936 20852 12000
rect 20916 11936 20932 12000
rect 20996 11936 21012 12000
rect 21076 11936 21092 12000
rect 21156 11936 21164 12000
rect 20844 10912 21164 11936
rect 20844 10848 20852 10912
rect 20916 10848 20932 10912
rect 20996 10848 21012 10912
rect 21076 10848 21092 10912
rect 21156 10848 21164 10912
rect 20844 9824 21164 10848
rect 20844 9760 20852 9824
rect 20916 9760 20932 9824
rect 20996 9760 21012 9824
rect 21076 9760 21092 9824
rect 21156 9760 21164 9824
rect 20844 8736 21164 9760
rect 20844 8672 20852 8736
rect 20916 8672 20932 8736
rect 20996 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21164 8736
rect 20844 7648 21164 8672
rect 20844 7584 20852 7648
rect 20916 7584 20932 7648
rect 20996 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21164 7648
rect 20844 6560 21164 7584
rect 20844 6496 20852 6560
rect 20916 6496 20932 6560
rect 20996 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21164 6560
rect 20844 5472 21164 6496
rect 20844 5408 20852 5472
rect 20916 5408 20932 5472
rect 20996 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21164 5472
rect 20844 4384 21164 5408
rect 20844 4320 20852 4384
rect 20916 4320 20932 4384
rect 20996 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21164 4384
rect 20844 3296 21164 4320
rect 20844 3232 20852 3296
rect 20916 3232 20932 3296
rect 20996 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21164 3296
rect 20844 2208 21164 3232
rect 20844 2144 20852 2208
rect 20916 2144 20932 2208
rect 20996 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21164 2208
rect 20844 2128 21164 2144
rect 22344 13632 22664 14656
rect 22344 13568 22352 13632
rect 22416 13568 22432 13632
rect 22496 13568 22512 13632
rect 22576 13568 22592 13632
rect 22656 13568 22664 13632
rect 22344 12544 22664 13568
rect 22344 12480 22352 12544
rect 22416 12480 22432 12544
rect 22496 12480 22512 12544
rect 22576 12480 22592 12544
rect 22656 12480 22664 12544
rect 22344 11456 22664 12480
rect 22344 11392 22352 11456
rect 22416 11392 22432 11456
rect 22496 11392 22512 11456
rect 22576 11392 22592 11456
rect 22656 11392 22664 11456
rect 22344 10368 22664 11392
rect 22344 10304 22352 10368
rect 22416 10304 22432 10368
rect 22496 10304 22512 10368
rect 22576 10304 22592 10368
rect 22656 10304 22664 10368
rect 22344 9280 22664 10304
rect 22344 9216 22352 9280
rect 22416 9216 22432 9280
rect 22496 9216 22512 9280
rect 22576 9216 22592 9280
rect 22656 9216 22664 9280
rect 22344 8192 22664 9216
rect 22344 8128 22352 8192
rect 22416 8128 22432 8192
rect 22496 8128 22512 8192
rect 22576 8128 22592 8192
rect 22656 8128 22664 8192
rect 22344 7104 22664 8128
rect 22344 7040 22352 7104
rect 22416 7040 22432 7104
rect 22496 7040 22512 7104
rect 22576 7040 22592 7104
rect 22656 7040 22664 7104
rect 22344 6016 22664 7040
rect 22344 5952 22352 6016
rect 22416 5952 22432 6016
rect 22496 5952 22512 6016
rect 22576 5952 22592 6016
rect 22656 5952 22664 6016
rect 22344 4928 22664 5952
rect 22344 4864 22352 4928
rect 22416 4864 22432 4928
rect 22496 4864 22512 4928
rect 22576 4864 22592 4928
rect 22656 4864 22664 4928
rect 22344 3840 22664 4864
rect 22344 3776 22352 3840
rect 22416 3776 22432 3840
rect 22496 3776 22512 3840
rect 22576 3776 22592 3840
rect 22656 3776 22664 3840
rect 22344 2752 22664 3776
rect 22344 2688 22352 2752
rect 22416 2688 22432 2752
rect 22496 2688 22512 2752
rect 22576 2688 22592 2752
rect 22656 2688 22664 2752
rect 22344 2128 22664 2688
rect 23844 25056 24164 25072
rect 23844 24992 23852 25056
rect 23916 24992 23932 25056
rect 23996 24992 24012 25056
rect 24076 24992 24092 25056
rect 24156 24992 24164 25056
rect 23844 23968 24164 24992
rect 23844 23904 23852 23968
rect 23916 23904 23932 23968
rect 23996 23904 24012 23968
rect 24076 23904 24092 23968
rect 24156 23904 24164 23968
rect 23844 22880 24164 23904
rect 23844 22816 23852 22880
rect 23916 22816 23932 22880
rect 23996 22816 24012 22880
rect 24076 22816 24092 22880
rect 24156 22816 24164 22880
rect 23844 21792 24164 22816
rect 23844 21728 23852 21792
rect 23916 21728 23932 21792
rect 23996 21728 24012 21792
rect 24076 21728 24092 21792
rect 24156 21728 24164 21792
rect 23844 20704 24164 21728
rect 23844 20640 23852 20704
rect 23916 20640 23932 20704
rect 23996 20640 24012 20704
rect 24076 20640 24092 20704
rect 24156 20640 24164 20704
rect 23844 19616 24164 20640
rect 23844 19552 23852 19616
rect 23916 19552 23932 19616
rect 23996 19552 24012 19616
rect 24076 19552 24092 19616
rect 24156 19552 24164 19616
rect 23844 18528 24164 19552
rect 23844 18464 23852 18528
rect 23916 18464 23932 18528
rect 23996 18464 24012 18528
rect 24076 18464 24092 18528
rect 24156 18464 24164 18528
rect 23844 17440 24164 18464
rect 23844 17376 23852 17440
rect 23916 17376 23932 17440
rect 23996 17376 24012 17440
rect 24076 17376 24092 17440
rect 24156 17376 24164 17440
rect 23844 16352 24164 17376
rect 23844 16288 23852 16352
rect 23916 16288 23932 16352
rect 23996 16288 24012 16352
rect 24076 16288 24092 16352
rect 24156 16288 24164 16352
rect 23844 15264 24164 16288
rect 23844 15200 23852 15264
rect 23916 15200 23932 15264
rect 23996 15200 24012 15264
rect 24076 15200 24092 15264
rect 24156 15200 24164 15264
rect 23844 14176 24164 15200
rect 23844 14112 23852 14176
rect 23916 14112 23932 14176
rect 23996 14112 24012 14176
rect 24076 14112 24092 14176
rect 24156 14112 24164 14176
rect 23844 13088 24164 14112
rect 23844 13024 23852 13088
rect 23916 13024 23932 13088
rect 23996 13024 24012 13088
rect 24076 13024 24092 13088
rect 24156 13024 24164 13088
rect 23844 12000 24164 13024
rect 23844 11936 23852 12000
rect 23916 11936 23932 12000
rect 23996 11936 24012 12000
rect 24076 11936 24092 12000
rect 24156 11936 24164 12000
rect 23844 10912 24164 11936
rect 23844 10848 23852 10912
rect 23916 10848 23932 10912
rect 23996 10848 24012 10912
rect 24076 10848 24092 10912
rect 24156 10848 24164 10912
rect 23844 9824 24164 10848
rect 23844 9760 23852 9824
rect 23916 9760 23932 9824
rect 23996 9760 24012 9824
rect 24076 9760 24092 9824
rect 24156 9760 24164 9824
rect 23844 8736 24164 9760
rect 23844 8672 23852 8736
rect 23916 8672 23932 8736
rect 23996 8672 24012 8736
rect 24076 8672 24092 8736
rect 24156 8672 24164 8736
rect 23844 7648 24164 8672
rect 23844 7584 23852 7648
rect 23916 7584 23932 7648
rect 23996 7584 24012 7648
rect 24076 7584 24092 7648
rect 24156 7584 24164 7648
rect 23844 6560 24164 7584
rect 23844 6496 23852 6560
rect 23916 6496 23932 6560
rect 23996 6496 24012 6560
rect 24076 6496 24092 6560
rect 24156 6496 24164 6560
rect 23844 5472 24164 6496
rect 23844 5408 23852 5472
rect 23916 5408 23932 5472
rect 23996 5408 24012 5472
rect 24076 5408 24092 5472
rect 24156 5408 24164 5472
rect 23844 4384 24164 5408
rect 23844 4320 23852 4384
rect 23916 4320 23932 4384
rect 23996 4320 24012 4384
rect 24076 4320 24092 4384
rect 24156 4320 24164 4384
rect 23844 3296 24164 4320
rect 23844 3232 23852 3296
rect 23916 3232 23932 3296
rect 23996 3232 24012 3296
rect 24076 3232 24092 3296
rect 24156 3232 24164 3296
rect 23844 2208 24164 3232
rect 23844 2144 23852 2208
rect 23916 2144 23932 2208
rect 23996 2144 24012 2208
rect 24076 2144 24092 2208
rect 24156 2144 24164 2208
rect 23844 2128 24164 2144
use sky130_fd_sc_hd__clkbuf_2  _389_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _391_
timestamp 1704896540
transform 1 0 12696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _392_
timestamp 1704896540
transform -1 0 10120 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _394_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _395_
timestamp 1704896540
transform -1 0 8924 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp 1704896540
transform 1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _397_
timestamp 1704896540
transform -1 0 5612 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1704896540
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _399_
timestamp 1704896540
transform 1 0 3312 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1704896540
transform 1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _401_
timestamp 1704896540
transform 1 0 7360 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1704896540
transform 1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _403_
timestamp 1704896540
transform -1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _404_
timestamp 1704896540
transform -1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _405_
timestamp 1704896540
transform -1 0 6532 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1704896540
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _407_
timestamp 1704896540
transform -1 0 11224 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp 1704896540
transform 1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _409_
timestamp 1704896540
transform -1 0 7084 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1704896540
transform 1 0 7820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _411_
timestamp 1704896540
transform -1 0 7084 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _412_
timestamp 1704896540
transform -1 0 7452 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _413_
timestamp 1704896540
transform -1 0 7084 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _414_
timestamp 1704896540
transform 1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _415_
timestamp 1704896540
transform -1 0 11040 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1704896540
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _417_
timestamp 1704896540
transform -1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _418_
timestamp 1704896540
transform -1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _419_
timestamp 1704896540
transform -1 0 11960 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1704896540
transform -1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _421_
timestamp 1704896540
transform -1 0 15548 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1704896540
transform 1 0 15180 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _423_
timestamp 1704896540
transform 1 0 14076 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1704896540
transform -1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _425_
timestamp 1704896540
transform -1 0 19872 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1704896540
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _427_
timestamp 1704896540
transform -1 0 15824 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1704896540
transform 1 0 16192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _429_
timestamp 1704896540
transform -1 0 20056 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _430_
timestamp 1704896540
transform -1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _431_
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _432_
timestamp 1704896540
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _433_
timestamp 1704896540
transform -1 0 19780 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1704896540
transform -1 0 20056 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _435_
timestamp 1704896540
transform -1 0 18584 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _436_
timestamp 1704896540
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _437_
timestamp 1704896540
transform -1 0 23736 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1704896540
transform -1 0 22172 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _439_
timestamp 1704896540
transform -1 0 23000 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1704896540
transform -1 0 22172 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _441_
timestamp 1704896540
transform -1 0 23736 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1704896540
transform -1 0 23184 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _443_
timestamp 1704896540
transform -1 0 18492 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1704896540
transform -1 0 18768 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _445_
timestamp 1704896540
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _446_
timestamp 1704896540
transform -1 0 16284 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _447_
timestamp 1704896540
transform -1 0 22632 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1704896540
transform -1 0 22908 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _449_
timestamp 1704896540
transform -1 0 19504 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _450_
timestamp 1704896540
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _451_
timestamp 1704896540
transform -1 0 17572 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _452_
timestamp 1704896540
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _453_
timestamp 1704896540
transform 1 0 19320 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _454_
timestamp 1704896540
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _455_
timestamp 1704896540
transform -1 0 17204 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _456_
timestamp 1704896540
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _457_
timestamp 1704896540
transform 1 0 19780 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _458_
timestamp 1704896540
transform -1 0 21712 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _459_
timestamp 1704896540
transform -1 0 16008 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _460_
timestamp 1704896540
transform -1 0 15088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _461_
timestamp 1704896540
transform -1 0 13984 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _462_
timestamp 1704896540
transform -1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _463_
timestamp 1704896540
transform -1 0 12512 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _464_
timestamp 1704896540
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13248 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _466_
timestamp 1704896540
transform -1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _467_
timestamp 1704896540
transform -1 0 8648 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1704896540
transform 1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp 1704896540
transform 1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp 1704896540
transform -1 0 3404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp 1704896540
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp 1704896540
transform 1 0 2392 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _475_
timestamp 1704896540
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp 1704896540
transform 1 0 7360 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _477_
timestamp 1704896540
transform -1 0 6256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _478_
timestamp 1704896540
transform 1 0 3956 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _479_
timestamp 1704896540
transform 1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _480_
timestamp 1704896540
transform -1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1704896540
transform 1 0 8924 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1704896540
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp 1704896540
transform 1 0 4232 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _484_
timestamp 1704896540
transform -1 0 3496 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 1704896540
transform 1 0 4692 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _486_
timestamp 1704896540
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _487_
timestamp 1704896540
transform 1 0 4140 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _488_
timestamp 1704896540
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _489_
timestamp 1704896540
transform 1 0 8280 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _490_
timestamp 1704896540
transform 1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 1704896540
transform 1 0 8924 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _492_
timestamp 1704896540
transform 1 0 8280 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _493_
timestamp 1704896540
transform 1 0 14168 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _494_
timestamp 1704896540
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _495_
timestamp 1704896540
transform 1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _496_
timestamp 1704896540
transform 1 0 13984 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _497_
timestamp 1704896540
transform 1 0 12420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _498_
timestamp 1704896540
transform 1 0 17112 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp 1704896540
transform 1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _500_
timestamp 1704896540
transform 1 0 13064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _501_
timestamp 1704896540
transform -1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _502_
timestamp 1704896540
transform 1 0 17204 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _503_
timestamp 1704896540
transform -1 0 16560 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _504_
timestamp 1704896540
transform 1 0 17756 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _505_
timestamp 1704896540
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _506_
timestamp 1704896540
transform 1 0 14168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _507_
timestamp 1704896540
transform 1 0 16008 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _508_
timestamp 1704896540
transform -1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _509_
timestamp 1704896540
transform 1 0 19872 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _510_
timestamp 1704896540
transform -1 0 19136 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _511_
timestamp 1704896540
transform 1 0 20792 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _512_
timestamp 1704896540
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _513_
timestamp 1704896540
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _514_
timestamp 1704896540
transform 1 0 20240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _515_
timestamp 1704896540
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _516_
timestamp 1704896540
transform 1 0 15180 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _517_
timestamp 1704896540
transform 1 0 20884 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _518_
timestamp 1704896540
transform 1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _519_
timestamp 1704896540
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _520_
timestamp 1704896540
transform 1 0 17572 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1704896540
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1704896540
transform 1 0 14628 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1704896540
transform -1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 1704896540
transform 1 0 19228 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1704896540
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _526_
timestamp 1704896540
transform 1 0 14904 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1704896540
transform 1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _528_
timestamp 1704896540
transform 1 0 18676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _529_
timestamp 1704896540
transform -1 0 19044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _530_
timestamp 1704896540
transform 1 0 13156 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _531_
timestamp 1704896540
transform -1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _532_
timestamp 1704896540
transform 1 0 10488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _533_
timestamp 1704896540
transform 1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _534_
timestamp 1704896540
transform 1 0 9936 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _535_
timestamp 1704896540
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _536_
timestamp 1704896540
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _537_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12512 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  _538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _539_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12696 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _540_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12052 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1704896540
transform -1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _542_
timestamp 1704896540
transform 1 0 12696 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _543_
timestamp 1704896540
transform -1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _544_
timestamp 1704896540
transform -1 0 10764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _546_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _548_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13248 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _549_
timestamp 1704896540
transform -1 0 14444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _550_
timestamp 1704896540
transform -1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1704896540
transform 1 0 4692 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1704896540
transform -1 0 3680 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1704896540
transform 1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1704896540
transform -1 0 7360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1704896540
transform 1 0 4600 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1704896540
transform -1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1704896540
transform 1 0 4048 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1704896540
transform -1 0 3312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1704896540
transform -1 0 9752 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1704896540
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _561_
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1704896540
transform 1 0 5060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _563_
timestamp 1704896540
transform -1 0 11408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _564_
timestamp 1704896540
transform 1 0 10120 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1704896540
transform -1 0 9936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _566_
timestamp 1704896540
transform -1 0 6256 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1704896540
transform -1 0 7360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _568_
timestamp 1704896540
transform -1 0 7176 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1704896540
transform -1 0 8004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _570_
timestamp 1704896540
transform -1 0 7268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1704896540
transform -1 0 7360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _572_
timestamp 1704896540
transform 1 0 9844 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1704896540
transform -1 0 9568 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _574_
timestamp 1704896540
transform 1 0 10212 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1704896540
transform -1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _576_
timestamp 1704896540
transform -1 0 16376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _577_
timestamp 1704896540
transform 1 0 15548 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1704896540
transform 1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _579_
timestamp 1704896540
transform -1 0 16192 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _580_
timestamp 1704896540
transform -1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _581_
timestamp 1704896540
transform -1 0 19136 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _582_
timestamp 1704896540
transform -1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _583_
timestamp 1704896540
transform -1 0 16376 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1704896540
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _585_
timestamp 1704896540
transform 1 0 20700 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _586_
timestamp 1704896540
transform 1 0 20056 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _587_
timestamp 1704896540
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1704896540
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _589_
timestamp 1704896540
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _590_
timestamp 1704896540
transform 1 0 17204 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _591_
timestamp 1704896540
transform 1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _592_
timestamp 1704896540
transform -1 0 21896 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _593_
timestamp 1704896540
transform -1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _594_
timestamp 1704896540
transform 1 0 22816 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _595_
timestamp 1704896540
transform -1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _596_
timestamp 1704896540
transform -1 0 22908 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _597_
timestamp 1704896540
transform 1 0 23184 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _598_
timestamp 1704896540
transform 1 0 18400 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _599_
timestamp 1704896540
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _600_
timestamp 1704896540
transform 1 0 21988 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _601_
timestamp 1704896540
transform -1 0 21712 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _602_
timestamp 1704896540
transform 1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _603_
timestamp 1704896540
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _604_
timestamp 1704896540
transform -1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _605_
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _606_
timestamp 1704896540
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _607_
timestamp 1704896540
transform -1 0 20884 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _608_
timestamp 1704896540
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _609_
timestamp 1704896540
transform -1 0 17480 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _610_
timestamp 1704896540
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _611_
timestamp 1704896540
transform 1 0 20792 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _612_
timestamp 1704896540
transform -1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _613_
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _614_
timestamp 1704896540
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _615_
timestamp 1704896540
transform 1 0 13984 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _616_
timestamp 1704896540
transform 1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _617_
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _618_
timestamp 1704896540
transform -1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _619_
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _620_
timestamp 1704896540
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _621_
timestamp 1704896540
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _622_
timestamp 1704896540
transform -1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _623_
timestamp 1704896540
transform 1 0 5796 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _624_
timestamp 1704896540
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _625_
timestamp 1704896540
transform 1 0 3680 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _626_
timestamp 1704896540
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _627_
timestamp 1704896540
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _628_
timestamp 1704896540
transform -1 0 7268 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _629_
timestamp 1704896540
transform -1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _630_
timestamp 1704896540
transform 1 0 5336 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _631_
timestamp 1704896540
transform 1 0 5244 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _632_
timestamp 1704896540
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _633_
timestamp 1704896540
transform 1 0 10488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _634_
timestamp 1704896540
transform 1 0 6348 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _635_
timestamp 1704896540
transform -1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _636_
timestamp 1704896540
transform 1 0 6348 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _637_
timestamp 1704896540
transform 1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _638_
timestamp 1704896540
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _639_
timestamp 1704896540
transform 1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _640_
timestamp 1704896540
transform 1 0 11040 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _641_
timestamp 1704896540
transform 1 0 10212 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _642_
timestamp 1704896540
transform -1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _643_
timestamp 1704896540
transform 1 0 10488 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _644_
timestamp 1704896540
transform -1 0 9936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _645_
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _646_
timestamp 1704896540
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _647_
timestamp 1704896540
transform 1 0 14352 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _648_
timestamp 1704896540
transform -1 0 13984 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _649_
timestamp 1704896540
transform 1 0 19872 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _650_
timestamp 1704896540
transform -1 0 19044 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _651_
timestamp 1704896540
transform 1 0 14260 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _652_
timestamp 1704896540
transform -1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _653_
timestamp 1704896540
transform -1 0 19136 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _654_
timestamp 1704896540
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _655_
timestamp 1704896540
transform 1 0 16744 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _656_
timestamp 1704896540
transform -1 0 19044 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _657_
timestamp 1704896540
transform 1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _658_
timestamp 1704896540
transform 1 0 18308 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _659_
timestamp 1704896540
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _660_
timestamp 1704896540
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _661_
timestamp 1704896540
transform -1 0 21712 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _662_
timestamp 1704896540
transform -1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _663_
timestamp 1704896540
transform 1 0 23368 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _664_
timestamp 1704896540
transform -1 0 22632 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _665_
timestamp 1704896540
transform 1 0 22632 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _666_
timestamp 1704896540
transform 1 0 17204 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _667_
timestamp 1704896540
transform -1 0 16560 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _668_
timestamp 1704896540
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _669_
timestamp 1704896540
transform 1 0 21804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 1704896540
transform 1 0 21068 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _671_
timestamp 1704896540
transform 1 0 18400 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp 1704896540
transform -1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _673_
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _674_
timestamp 1704896540
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _675_
timestamp 1704896540
transform -1 0 20516 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _676_
timestamp 1704896540
transform 1 0 21620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _677_
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _678_
timestamp 1704896540
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _679_
timestamp 1704896540
transform -1 0 21160 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _680_
timestamp 1704896540
transform -1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _681_
timestamp 1704896540
transform 1 0 14260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _682_
timestamp 1704896540
transform 1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _683_
timestamp 1704896540
transform 1 0 12604 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _684_
timestamp 1704896540
transform -1 0 12052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _685_
timestamp 1704896540
transform 1 0 10580 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _686_
timestamp 1704896540
transform -1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _687_
timestamp 1704896540
transform 1 0 12696 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _688_
timestamp 1704896540
transform -1 0 13984 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _689_
timestamp 1704896540
transform -1 0 8280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _690_
timestamp 1704896540
transform 1 0 2392 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _691_
timestamp 1704896540
transform 1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _692_
timestamp 1704896540
transform -1 0 6256 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1704896540
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _694_
timestamp 1704896540
transform 1 0 2668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _695_
timestamp 1704896540
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _696_
timestamp 1704896540
transform 1 0 2392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _697_
timestamp 1704896540
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _698_
timestamp 1704896540
transform 1 0 6532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _699_
timestamp 1704896540
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _700_
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _701_
timestamp 1704896540
transform -1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _702_
timestamp 1704896540
transform -1 0 8372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _703_
timestamp 1704896540
transform 1 0 8924 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _704_
timestamp 1704896540
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _705_
timestamp 1704896540
transform 1 0 4324 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _706_
timestamp 1704896540
transform 1 0 3864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _707_
timestamp 1704896540
transform 1 0 4140 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _708_
timestamp 1704896540
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _709_
timestamp 1704896540
transform 1 0 4600 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _710_
timestamp 1704896540
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _711_
timestamp 1704896540
transform 1 0 8372 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _712_
timestamp 1704896540
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _713_
timestamp 1704896540
transform 1 0 8924 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _714_
timestamp 1704896540
transform 1 0 8280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _715_
timestamp 1704896540
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _716_
timestamp 1704896540
transform 1 0 12972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _717_
timestamp 1704896540
transform -1 0 12052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _718_
timestamp 1704896540
transform 1 0 13156 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _719_
timestamp 1704896540
transform 1 0 12696 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _720_
timestamp 1704896540
transform 1 0 17940 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _721_
timestamp 1704896540
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _722_
timestamp 1704896540
transform 1 0 13156 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _723_
timestamp 1704896540
transform 1 0 12696 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _724_
timestamp 1704896540
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _725_
timestamp 1704896540
transform -1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _726_
timestamp 1704896540
transform 1 0 17204 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _727_
timestamp 1704896540
transform 1 0 16744 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _728_
timestamp 1704896540
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _729_
timestamp 1704896540
transform 1 0 15364 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _730_
timestamp 1704896540
transform 1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _731_
timestamp 1704896540
transform 1 0 20608 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _732_
timestamp 1704896540
transform 1 0 19504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _733_
timestamp 1704896540
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _734_
timestamp 1704896540
transform 1 0 19780 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _735_
timestamp 1704896540
transform 1 0 20700 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _736_
timestamp 1704896540
transform 1 0 20516 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _737_
timestamp 1704896540
transform 1 0 15548 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _738_
timestamp 1704896540
transform 1 0 15180 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _739_
timestamp 1704896540
transform 1 0 21160 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _740_
timestamp 1704896540
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _741_
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _742_
timestamp 1704896540
transform 1 0 16744 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _743_
timestamp 1704896540
transform -1 0 16560 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _744_
timestamp 1704896540
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _745_
timestamp 1704896540
transform -1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _746_
timestamp 1704896540
transform -1 0 19136 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _747_
timestamp 1704896540
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _748_
timestamp 1704896540
transform 1 0 14168 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _749_
timestamp 1704896540
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _750_
timestamp 1704896540
transform 1 0 18308 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _751_
timestamp 1704896540
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _752_
timestamp 1704896540
transform 1 0 15364 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _753_
timestamp 1704896540
transform -1 0 12880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _754_
timestamp 1704896540
transform 1 0 11316 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _755_
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _756_
timestamp 1704896540
transform 1 0 9844 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp 1704896540
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _758_
timestamp 1704896540
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _759_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9292 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _761_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _762_
timestamp 1704896540
transform -1 0 8740 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _763_
timestamp 1704896540
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _764_
timestamp 1704896540
transform 1 0 8372 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _765_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _767_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _768_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _769_
timestamp 1704896540
transform 1 0 9476 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _770_
timestamp 1704896540
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _771_
timestamp 1704896540
transform 1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _772_
timestamp 1704896540
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _773_
timestamp 1704896540
transform 1 0 8004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _774_
timestamp 1704896540
transform 1 0 8372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _775_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _776_
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _777_
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _778_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand4bb_1  _779_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _780_
timestamp 1704896540
transform 1 0 6624 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _781_
timestamp 1704896540
transform -1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _782_
timestamp 1704896540
transform -1 0 6164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _783_
timestamp 1704896540
transform 1 0 5888 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _784_
timestamp 1704896540
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _785_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7912 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _786_
timestamp 1704896540
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _788_
timestamp 1704896540
transform 1 0 7728 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _789_
timestamp 1704896540
transform -1 0 7728 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _790_
timestamp 1704896540
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _792_
timestamp 1704896540
transform -1 0 11040 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _793_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7912 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _794_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _795_
timestamp 1704896540
transform -1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _796_
timestamp 1704896540
transform -1 0 10948 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _797_
timestamp 1704896540
transform -1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _798_
timestamp 1704896540
transform -1 0 11592 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _799_
timestamp 1704896540
transform 1 0 10028 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _800_
timestamp 1704896540
transform 1 0 9476 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _801_
timestamp 1704896540
transform 1 0 9844 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _803_
timestamp 1704896540
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _805_
timestamp 1704896540
transform 1 0 8648 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _806_
timestamp 1704896540
transform 1 0 9292 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _807_
timestamp 1704896540
transform -1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _809_
timestamp 1704896540
transform 1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1472 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1704896540
transform 1 0 5428 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1704896540
transform 1 0 1840 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1704896540
transform 1 0 1472 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1704896540
transform 1 0 2484 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1704896540
transform 1 0 7912 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1704896540
transform 1 0 3772 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1704896540
transform 1 0 3220 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp 1704896540
transform 1 0 3128 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp 1704896540
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp 1704896540
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp 1704896540
transform 1 0 12052 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp 1704896540
transform 1 0 12236 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp 1704896540
transform 1 0 16468 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp 1704896540
transform 1 0 12144 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp 1704896540
transform 1 0 16652 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp 1704896540
transform 1 0 16284 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp 1704896540
transform 1 0 14536 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp 1704896540
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp 1704896540
transform 1 0 19320 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp 1704896540
transform 1 0 20056 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp 1704896540
transform 1 0 14812 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _833_
timestamp 1704896540
transform 1 0 19412 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _834_
timestamp 1704896540
transform 1 0 16008 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _836_
timestamp 1704896540
transform 1 0 17756 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp 1704896540
transform 1 0 13432 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _838_
timestamp 1704896540
transform 1 0 19688 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp 1704896540
transform 1 0 12512 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp 1704896540
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _841_
timestamp 1704896540
transform 1 0 9108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _843_
timestamp 1704896540
transform 1 0 10120 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _844_
timestamp 1704896540
transform 1 0 3956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _845_
timestamp 1704896540
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _846_
timestamp 1704896540
transform 1 0 4324 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _847_
timestamp 1704896540
transform -1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _848_
timestamp 1704896540
transform -1 0 9568 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _849_
timestamp 1704896540
transform 1 0 4784 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _850_
timestamp 1704896540
transform 1 0 9936 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _851_
timestamp 1704896540
transform -1 0 7820 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _852_
timestamp 1704896540
transform -1 0 8556 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _853_
timestamp 1704896540
transform -1 0 8556 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _854_
timestamp 1704896540
transform 1 0 9568 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _855_
timestamp 1704896540
transform 1 0 9936 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _856_
timestamp 1704896540
transform 1 0 14536 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _857_
timestamp 1704896540
transform -1 0 16468 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp 1704896540
transform -1 0 20700 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp 1704896540
transform -1 0 16192 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp 1704896540
transform 1 0 19136 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp 1704896540
transform -1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp 1704896540
transform 1 0 17112 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp 1704896540
transform 1 0 21896 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp 1704896540
transform 1 0 21896 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp 1704896540
transform 1 0 22172 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1704896540
transform 1 0 17296 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp 1704896540
transform 1 0 22172 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp 1704896540
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp 1704896540
transform 1 0 16008 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp 1704896540
transform -1 0 21436 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp 1704896540
transform 1 0 15640 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp 1704896540
transform 1 0 21712 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp 1704896540
transform 1 0 14168 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp 1704896540
transform 1 0 12512 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp 1704896540
transform -1 0 12972 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp 1704896540
transform 1 0 3220 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp 1704896540
transform 1 0 6900 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp 1704896540
transform 1 0 3956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp 1704896540
transform -1 0 8740 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp 1704896540
transform 1 0 4784 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp 1704896540
transform 1 0 9936 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp 1704896540
transform 1 0 5612 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp 1704896540
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp 1704896540
transform 1 0 5336 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp 1704896540
transform 1 0 9936 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 1704896540
transform 1 0 9936 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 1704896540
transform 1 0 13248 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 1704896540
transform 1 0 13892 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 1704896540
transform 1 0 19228 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 1704896540
transform 1 0 14076 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 1704896540
transform 1 0 19228 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 1704896540
transform 1 0 18032 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 1704896540
transform 1 0 16836 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp 1704896540
transform 1 0 21804 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp 1704896540
transform -1 0 23276 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 1704896540
transform 1 0 21712 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 1704896540
transform 1 0 16928 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 1704896540
transform 1 0 20884 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 1704896540
transform 1 0 17480 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1704896540
transform -1 0 18124 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1704896540
transform -1 0 20884 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 1704896540
transform -1 0 18676 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 1704896540
transform -1 0 21712 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 1704896540
transform 1 0 12788 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 1704896540
transform 1 0 12328 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 1704896540
transform -1 0 13984 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 1704896540
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 1704896540
transform -1 0 7084 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 1704896540
transform 1 0 1840 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 1704896540
transform 1 0 1472 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 1704896540
transform 1 0 5888 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 1704896540
transform 1 0 2208 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 1704896540
transform 1 0 8004 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _915_
timestamp 1704896540
transform 1 0 3496 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _916_
timestamp 1704896540
transform 1 0 3220 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _917_
timestamp 1704896540
transform 1 0 3220 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _918_
timestamp 1704896540
transform 1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _919_
timestamp 1704896540
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _920_
timestamp 1704896540
transform 1 0 12052 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _921_
timestamp 1704896540
transform 1 0 12236 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _922_
timestamp 1704896540
transform 1 0 16468 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _923_
timestamp 1704896540
transform 1 0 12236 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _924_
timestamp 1704896540
transform 1 0 16744 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _925_
timestamp 1704896540
transform 1 0 16376 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 1704896540
transform 1 0 14536 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 1704896540
transform 1 0 19136 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 1704896540
transform 1 0 19320 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 1704896540
transform 1 0 20148 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 1704896540
transform 1 0 14812 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 1704896540
transform 1 0 19688 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _932_
timestamp 1704896540
transform 1 0 16376 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 1704896540
transform 1 0 14076 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 1704896540
transform 1 0 13432 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 1704896540
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 1704896540
transform 1 0 12880 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _938_
timestamp 1704896540
transform 1 0 10580 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _939_
timestamp 1704896540
transform 1 0 9108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _940_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6440 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _941_
timestamp 1704896540
transform 1 0 9476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _942_
timestamp 1704896540
transform 1 0 6072 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _943_
timestamp 1704896540
transform 1 0 4692 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _944_
timestamp 1704896540
transform 1 0 5244 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _945_
timestamp 1704896540
transform 1 0 6624 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _946_
timestamp 1704896540
transform -1 0 13340 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _947_
timestamp 1704896540
transform -1 0 13524 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _948_
timestamp 1704896540
transform 1 0 10488 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _949_
timestamp 1704896540
transform 1 0 10212 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_Clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12512 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_Clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6256 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_Clk
timestamp 1704896540
transform -1 0 3956 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_Clk
timestamp 1704896540
transform 1 0 8188 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_Clk
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_Clk
timestamp 1704896540
transform 1 0 5152 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_Clk
timestamp 1704896540
transform -1 0 7728 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_Clk
timestamp 1704896540
transform 1 0 10764 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_Clk
timestamp 1704896540
transform 1 0 11224 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_Clk
timestamp 1704896540
transform -1 0 15272 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_Clk
timestamp 1704896540
transform 1 0 14352 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_Clk
timestamp 1704896540
transform -1 0 20792 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_Clk
timestamp 1704896540
transform -1 0 20516 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_Clk
timestamp 1704896540
transform 1 0 16652 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_Clk
timestamp 1704896540
transform 1 0 16836 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_Clk
timestamp 1704896540
transform 1 0 21804 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_Clk
timestamp 1704896540
transform 1 0 20700 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  clkload0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  clkload1
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinvlp_2  clkload2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  clkload3
timestamp 1704896540
transform -1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  clkload4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  clkload5
timestamp 1704896540
transform -1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 1704896540
transform -1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_2  clkload7
timestamp 1704896540
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15088 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload9
timestamp 1704896540
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload10
timestamp 1704896540
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload11
timestamp 1704896540
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload12
timestamp 1704896540
transform -1 0 17204 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload13
timestamp 1704896540
transform -1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20700 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 1704896540
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout75
timestamp 1704896540
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1704896540
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_118 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_128
timestamp 1704896540
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_146
timestamp 1704896540
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_156
timestamp 1704896540
transform 1 0 15456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_160
timestamp 1704896540
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1704896540
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1704896540
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_184
timestamp 1704896540
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_188
timestamp 1704896540
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_202
timestamp 1704896540
transform 1 0 19688 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_214
timestamp 1704896540
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1704896540
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_231
timestamp 1704896540
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_243
timestamp 1704896540
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_80
timestamp 1704896540
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_95
timestamp 1704896540
transform 1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_116
timestamp 1704896540
transform 1 0 11776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_128 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12880 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_162
timestamp 1704896540
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_215
timestamp 1704896540
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_237
timestamp 1704896540
transform 1 0 22908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_245
timestamp 1704896540
transform 1 0 23644 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_72
timestamp 1704896540
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_114
timestamp 1704896540
transform 1 0 11592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_135
timestamp 1704896540
transform 1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1704896540
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_229
timestamp 1704896540
transform 1 0 22172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_241
timestamp 1704896540
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_245
timestamp 1704896540
transform 1 0 23644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_47
timestamp 1704896540
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_60
timestamp 1704896540
transform 1 0 6624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_68
timestamp 1704896540
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_74
timestamp 1704896540
transform 1 0 7912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_91
timestamp 1704896540
transform 1 0 9476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_133
timestamp 1704896540
transform 1 0 13340 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1704896540
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_197
timestamp 1704896540
transform 1 0 19228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1704896540
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_233
timestamp 1704896540
transform 1 0 22540 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_245
timestamp 1704896540
transform 1 0 23644 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_49
timestamp 1704896540
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_61
timestamp 1704896540
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1704896540
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_100
timestamp 1704896540
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_108
timestamp 1704896540
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_120
timestamp 1704896540
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 1704896540
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1704896540
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1704896540
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_182
timestamp 1704896540
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_186
timestamp 1704896540
transform 1 0 18216 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1704896540
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1704896540
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_245
timestamp 1704896540
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_47
timestamp 1704896540
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_68
timestamp 1704896540
transform 1 0 7360 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_89
timestamp 1704896540
transform 1 0 9292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_101
timestamp 1704896540
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1704896540
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_153
timestamp 1704896540
transform 1 0 15180 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_162
timestamp 1704896540
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_186
timestamp 1704896540
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_198
timestamp 1704896540
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_219
timestamp 1704896540
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_245
timestamp 1704896540
transform 1 0 23644 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1704896540
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_95
timestamp 1704896540
transform 1 0 9844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_99
timestamp 1704896540
transform 1 0 10212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_111
timestamp 1704896540
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1704896540
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1704896540
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1704896540
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_179
timestamp 1704896540
transform 1 0 17572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_187
timestamp 1704896540
transform 1 0 18308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_223
timestamp 1704896540
transform 1 0 21620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_235
timestamp 1704896540
transform 1 0 22724 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_243
timestamp 1704896540
transform 1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_75
timestamp 1704896540
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_89
timestamp 1704896540
transform 1 0 9292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_133
timestamp 1704896540
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1704896540
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 1704896540
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_37
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_49
timestamp 1704896540
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_89
timestamp 1704896540
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_96
timestamp 1704896540
transform 1 0 9936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_100
timestamp 1704896540
transform 1 0 10304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_108
timestamp 1704896540
transform 1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_124
timestamp 1704896540
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_131
timestamp 1704896540
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_156
timestamp 1704896540
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_186
timestamp 1704896540
transform 1 0 18216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_240
timestamp 1704896540
transform 1 0 23184 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_25
timestamp 1704896540
transform 1 0 3404 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_47
timestamp 1704896540
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_90
timestamp 1704896540
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 1704896540
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1704896540
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1704896540
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_121
timestamp 1704896540
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_154
timestamp 1704896540
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_158
timestamp 1704896540
transform 1 0 15640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_189
timestamp 1704896540
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_233
timestamp 1704896540
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_241
timestamp 1704896540
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 1704896540
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_24
timestamp 1704896540
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_75
timestamp 1704896540
transform 1 0 8004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_131
timestamp 1704896540
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_135
timestamp 1704896540
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_149
timestamp 1704896540
transform 1 0 14812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_161
timestamp 1704896540
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_173
timestamp 1704896540
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_177
timestamp 1704896540
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1704896540
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1704896540
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_226
timestamp 1704896540
transform 1 0 21896 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_238
timestamp 1704896540
transform 1 0 23000 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_7
timestamp 1704896540
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1704896540
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_65
timestamp 1704896540
transform 1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_76
timestamp 1704896540
transform 1 0 8096 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_87
timestamp 1704896540
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_94
timestamp 1704896540
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_102
timestamp 1704896540
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1704896540
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_155
timestamp 1704896540
transform 1 0 15364 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_163
timestamp 1704896540
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_219
timestamp 1704896540
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1704896540
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1704896540
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_237
timestamp 1704896540
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_245
timestamp 1704896540
transform 1 0 23644 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_6
timestamp 1704896540
transform 1 0 1656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_15
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1704896540
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_37
timestamp 1704896540
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_47
timestamp 1704896540
transform 1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_61
timestamp 1704896540
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_73
timestamp 1704896540
transform 1 0 7820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1704896540
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_100
timestamp 1704896540
transform 1 0 10304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_122
timestamp 1704896540
transform 1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1704896540
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_213
timestamp 1704896540
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_231
timestamp 1704896540
transform 1 0 22356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_237
timestamp 1704896540
transform 1 0 22908 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_6
timestamp 1704896540
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_12
timestamp 1704896540
transform 1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_31
timestamp 1704896540
transform 1 0 3956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_41
timestamp 1704896540
transform 1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_66
timestamp 1704896540
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_88
timestamp 1704896540
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_96
timestamp 1704896540
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_104
timestamp 1704896540
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1704896540
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_164
timestamp 1704896540
transform 1 0 16192 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_178
timestamp 1704896540
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_215
timestamp 1704896540
transform 1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_220
timestamp 1704896540
transform 1 0 21344 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_45
timestamp 1704896540
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_93
timestamp 1704896540
transform 1 0 9660 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_119
timestamp 1704896540
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_190
timestamp 1704896540
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1704896540
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_209
timestamp 1704896540
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_20
timestamp 1704896540
transform 1 0 2944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_60
timestamp 1704896540
transform 1 0 6624 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_98
timestamp 1704896540
transform 1 0 10120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1704896540
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12604 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_130
timestamp 1704896540
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_142
timestamp 1704896540
transform 1 0 14168 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_148
timestamp 1704896540
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_160
timestamp 1704896540
transform 1 0 15824 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1704896540
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_177
timestamp 1704896540
transform 1 0 17388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_189
timestamp 1704896540
transform 1 0 18492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_197
timestamp 1704896540
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21804 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_245
timestamp 1704896540
transform 1 0 23644 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_23
timestamp 1704896540
transform 1 0 3220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_45
timestamp 1704896540
transform 1 0 5244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_79
timestamp 1704896540
transform 1 0 8372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_113
timestamp 1704896540
transform 1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_124
timestamp 1704896540
transform 1 0 12512 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_128
timestamp 1704896540
transform 1 0 12880 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_145
timestamp 1704896540
transform 1 0 14444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_151
timestamp 1704896540
transform 1 0 14996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_156
timestamp 1704896540
transform 1 0 15456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_164
timestamp 1704896540
transform 1 0 16192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_169
timestamp 1704896540
transform 1 0 16652 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_184
timestamp 1704896540
transform 1 0 18032 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 1704896540
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1704896540
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1704896540
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_244
timestamp 1704896540
transform 1 0 23552 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_6
timestamp 1704896540
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_18
timestamp 1704896540
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 1704896540
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_61
timestamp 1704896540
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_70
timestamp 1704896540
transform 1 0 7544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_122
timestamp 1704896540
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_198
timestamp 1704896540
transform 1 0 19320 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_210
timestamp 1704896540
transform 1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_234
timestamp 1704896540
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_6
timestamp 1704896540
transform 1 0 1656 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_18
timestamp 1704896540
transform 1 0 2760 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_24
timestamp 1704896540
transform 1 0 3312 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_32
timestamp 1704896540
transform 1 0 4048 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_44
timestamp 1704896540
transform 1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_56
timestamp 1704896540
transform 1 0 6256 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_68
timestamp 1704896540
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_80
timestamp 1704896540
transform 1 0 8464 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_221
timestamp 1704896540
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_241
timestamp 1704896540
transform 1 0 23276 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1704896540
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_47
timestamp 1704896540
transform 1 0 5428 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_81
timestamp 1704896540
transform 1 0 8556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_86
timestamp 1704896540
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_90
timestamp 1704896540
transform 1 0 9384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_94
timestamp 1704896540
transform 1 0 9752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_132
timestamp 1704896540
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_140
timestamp 1704896540
transform 1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_162
timestamp 1704896540
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_50
timestamp 1704896540
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1704896540
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_97
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_105
timestamp 1704896540
transform 1 0 10764 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_112
timestamp 1704896540
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_124
timestamp 1704896540
transform 1 0 12512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1704896540
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_149
timestamp 1704896540
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_172
timestamp 1704896540
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_180
timestamp 1704896540
transform 1 0 17664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_192
timestamp 1704896540
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_197
timestamp 1704896540
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_203
timestamp 1704896540
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_213
timestamp 1704896540
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_21
timestamp 1704896540
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_92
timestamp 1704896540
transform 1 0 9568 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_100
timestamp 1704896540
transform 1 0 10304 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1704896540
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_121
timestamp 1704896540
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_152
timestamp 1704896540
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_156
timestamp 1704896540
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_173
timestamp 1704896540
transform 1 0 17020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_185
timestamp 1704896540
transform 1 0 18124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_197
timestamp 1704896540
transform 1 0 19228 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_205
timestamp 1704896540
transform 1 0 19964 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1704896540
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 1704896540
transform 1 0 23644 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_7
timestamp 1704896540
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_12
timestamp 1704896540
transform 1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_23
timestamp 1704896540
transform 1 0 3220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_46
timestamp 1704896540
transform 1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_51
timestamp 1704896540
transform 1 0 5796 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_56
timestamp 1704896540
transform 1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_97
timestamp 1704896540
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_119
timestamp 1704896540
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_123
timestamp 1704896540
transform 1 0 12420 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_174
timestamp 1704896540
transform 1 0 17112 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_192
timestamp 1704896540
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_208
timestamp 1704896540
transform 1 0 20240 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_224
timestamp 1704896540
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_6
timestamp 1704896540
transform 1 0 1656 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_18
timestamp 1704896540
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_28
timestamp 1704896540
transform 1 0 3680 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_48
timestamp 1704896540
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_63
timestamp 1704896540
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1704896540
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_197
timestamp 1704896540
transform 1 0 19228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1704896540
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_241
timestamp 1704896540
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_6
timestamp 1704896540
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_18
timestamp 1704896540
transform 1 0 2760 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_22
timestamp 1704896540
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_38
timestamp 1704896540
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_56
timestamp 1704896540
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_68
timestamp 1704896540
transform 1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1704896540
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp 1704896540
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_101
timestamp 1704896540
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_120
timestamp 1704896540
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1704896540
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1704896540
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1704896540
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1704896540
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_6
timestamp 1704896540
transform 1 0 1656 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_78
timestamp 1704896540
transform 1 0 8280 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_90
timestamp 1704896540
transform 1 0 9384 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_102
timestamp 1704896540
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_131
timestamp 1704896540
transform 1 0 13156 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_143
timestamp 1704896540
transform 1 0 14260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_151
timestamp 1704896540
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1704896540
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_192
timestamp 1704896540
transform 1 0 18768 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_200
timestamp 1704896540
transform 1 0 19504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1704896540
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_245
timestamp 1704896540
transform 1 0 23644 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_7
timestamp 1704896540
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_11
timestamp 1704896540
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_62
timestamp 1704896540
transform 1 0 6808 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_91
timestamp 1704896540
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_96
timestamp 1704896540
transform 1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_102
timestamp 1704896540
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_108
timestamp 1704896540
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_112
timestamp 1704896540
transform 1 0 11408 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_117
timestamp 1704896540
transform 1 0 11868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_129
timestamp 1704896540
transform 1 0 12972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1704896540
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_150
timestamp 1704896540
transform 1 0 14904 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_162
timestamp 1704896540
transform 1 0 16008 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_171
timestamp 1704896540
transform 1 0 16836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_183
timestamp 1704896540
transform 1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1704896540
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1704896540
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_205
timestamp 1704896540
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_226
timestamp 1704896540
transform 1 0 21896 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_245
timestamp 1704896540
transform 1 0 23644 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_39
timestamp 1704896540
transform 1 0 4692 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1704896540
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_65
timestamp 1704896540
transform 1 0 7084 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_71
timestamp 1704896540
transform 1 0 7636 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_95
timestamp 1704896540
transform 1 0 9844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_131
timestamp 1704896540
transform 1 0 13156 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_160
timestamp 1704896540
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_173
timestamp 1704896540
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_211
timestamp 1704896540
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_225
timestamp 1704896540
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_245
timestamp 1704896540
transform 1 0 23644 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1704896540
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_41
timestamp 1704896540
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_45
timestamp 1704896540
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_62
timestamp 1704896540
transform 1 0 6808 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_117
timestamp 1704896540
transform 1 0 11868 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1704896540
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1704896540
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_162
timestamp 1704896540
transform 1 0 16008 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 1704896540
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_222
timestamp 1704896540
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_240
timestamp 1704896540
transform 1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_15
timestamp 1704896540
transform 1 0 2484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_21
timestamp 1704896540
transform 1 0 3036 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_47
timestamp 1704896540
transform 1 0 5428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1704896540
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1704896540
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_88
timestamp 1704896540
transform 1 0 9200 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_113
timestamp 1704896540
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_135
timestamp 1704896540
transform 1 0 13524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1704896540
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_180
timestamp 1704896540
transform 1 0 17664 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1704896540
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1704896540
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_18
timestamp 1704896540
transform 1 0 2760 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_24
timestamp 1704896540
transform 1 0 3312 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_32
timestamp 1704896540
transform 1 0 4048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_42
timestamp 1704896540
transform 1 0 4968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1704896540
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_93
timestamp 1704896540
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_104
timestamp 1704896540
transform 1 0 10672 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_116
timestamp 1704896540
transform 1 0 11776 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_127
timestamp 1704896540
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1704896540
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_152
timestamp 1704896540
transform 1 0 15088 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_182
timestamp 1704896540
transform 1 0 17848 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1704896540
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_206
timestamp 1704896540
transform 1 0 20056 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_223
timestamp 1704896540
transform 1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_7
timestamp 1704896540
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_19
timestamp 1704896540
transform 1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1704896540
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_77
timestamp 1704896540
transform 1 0 8188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_89
timestamp 1704896540
transform 1 0 9292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_98
timestamp 1704896540
transform 1 0 10120 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_116
timestamp 1704896540
transform 1 0 11776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_128
timestamp 1704896540
transform 1 0 12880 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_146
timestamp 1704896540
transform 1 0 14536 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_152
timestamp 1704896540
transform 1 0 15088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_156
timestamp 1704896540
transform 1 0 15456 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1704896540
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_172
timestamp 1704896540
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_180
timestamp 1704896540
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_189
timestamp 1704896540
transform 1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_197
timestamp 1704896540
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_208
timestamp 1704896540
transform 1 0 20240 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_214
timestamp 1704896540
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1704896540
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_241
timestamp 1704896540
transform 1 0 23276 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1704896540
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1704896540
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1704896540
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1704896540
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_65
timestamp 1704896540
transform 1 0 7084 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_69
timestamp 1704896540
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1704896540
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_94
timestamp 1704896540
transform 1 0 9752 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_107
timestamp 1704896540
transform 1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_120
timestamp 1704896540
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_132
timestamp 1704896540
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_141
timestamp 1704896540
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_164
timestamp 1704896540
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_168
timestamp 1704896540
transform 1 0 16560 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1704896540
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_200
timestamp 1704896540
transform 1 0 19504 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_212
timestamp 1704896540
transform 1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_224
timestamp 1704896540
transform 1 0 21712 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_232
timestamp 1704896540
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1704896540
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 1704896540
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_39
timestamp 1704896540
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_90
timestamp 1704896540
transform 1 0 9384 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_137
timestamp 1704896540
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_164
timestamp 1704896540
transform 1 0 16192 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_169
timestamp 1704896540
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_182
timestamp 1704896540
transform 1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_212
timestamp 1704896540
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1704896540
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_237
timestamp 1704896540
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_242
timestamp 1704896540
transform 1 0 23368 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1704896540
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_15
timestamp 1704896540
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_23
timestamp 1704896540
transform 1 0 3220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_32
timestamp 1704896540
transform 1 0 4048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_42
timestamp 1704896540
transform 1 0 4968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_88
timestamp 1704896540
transform 1 0 9200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_165
timestamp 1704896540
transform 1 0 16284 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1704896540
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_222
timestamp 1704896540
transform 1 0 21528 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_234
timestamp 1704896540
transform 1 0 22632 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1704896540
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_15
timestamp 1704896540
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_39
timestamp 1704896540
transform 1 0 4692 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1704896540
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_74
timestamp 1704896540
transform 1 0 7912 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_91
timestamp 1704896540
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_95
timestamp 1704896540
transform 1 0 9844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_130
timestamp 1704896540
transform 1 0 13064 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_149
timestamp 1704896540
transform 1 0 14812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1704896540
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1704896540
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_186
timestamp 1704896540
transform 1 0 18216 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_212
timestamp 1704896540
transform 1 0 20608 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1704896540
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1704896540
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_237
timestamp 1704896540
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_241
timestamp 1704896540
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1704896540
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1704896540
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1704896540
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 1704896540
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_56
timestamp 1704896540
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_75
timestamp 1704896540
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1704896540
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_105
timestamp 1704896540
transform 1 0 10764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_117
timestamp 1704896540
transform 1 0 11868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_129
timestamp 1704896540
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1704896540
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_157
timestamp 1704896540
transform 1 0 15548 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_171
timestamp 1704896540
transform 1 0 16836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_183
timestamp 1704896540
transform 1 0 17940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_187
timestamp 1704896540
transform 1 0 18308 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 1704896540
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 1704896540
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_210
timestamp 1704896540
transform 1 0 20424 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_222
timestamp 1704896540
transform 1 0 21528 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_234
timestamp 1704896540
transform 1 0 22632 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1704896540
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1704896540
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_27
timestamp 1704896540
transform 1 0 3588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_33
timestamp 1704896540
transform 1 0 4140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1704896540
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_66
timestamp 1704896540
transform 1 0 7176 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_98
timestamp 1704896540
transform 1 0 10120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1704896540
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1704896540
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_125
timestamp 1704896540
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_129
timestamp 1704896540
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_139
timestamp 1704896540
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_169
timestamp 1704896540
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_177
timestamp 1704896540
transform 1 0 17388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_189
timestamp 1704896540
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_196
timestamp 1704896540
transform 1 0 19136 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_208
timestamp 1704896540
transform 1 0 20240 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_220
timestamp 1704896540
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1704896540
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_237
timestamp 1704896540
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_245
timestamp 1704896540
transform 1 0 23644 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1704896540
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1704896540
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1704896540
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_29
timestamp 1704896540
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_33
timestamp 1704896540
transform 1 0 4140 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_76
timestamp 1704896540
transform 1 0 8096 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1704896540
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_94
timestamp 1704896540
transform 1 0 9752 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_118
timestamp 1704896540
transform 1 0 11960 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_136
timestamp 1704896540
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_166
timestamp 1704896540
transform 1 0 16376 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1704896540
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_213
timestamp 1704896540
transform 1 0 20700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_225
timestamp 1704896540
transform 1 0 21804 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_237
timestamp 1704896540
transform 1 0 22908 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_245
timestamp 1704896540
transform 1 0 23644 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1704896540
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_15
timestamp 1704896540
transform 1 0 2484 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_42
timestamp 1704896540
transform 1 0 4968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_73
timestamp 1704896540
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_137
timestamp 1704896540
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_172
timestamp 1704896540
transform 1 0 16928 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1704896540
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_237
timestamp 1704896540
transform 1 0 22908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_245
timestamp 1704896540
transform 1 0 23644 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1704896540
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1704896540
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1704896540
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_45
timestamp 1704896540
transform 1 0 5244 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_68
timestamp 1704896540
transform 1 0 7360 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_76
timestamp 1704896540
transform 1 0 8096 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_94
timestamp 1704896540
transform 1 0 9752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_124
timestamp 1704896540
transform 1 0 12512 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_129
timestamp 1704896540
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_141
timestamp 1704896540
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_183
timestamp 1704896540
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_213
timestamp 1704896540
transform 1 0 20700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_225
timestamp 1704896540
transform 1 0 21804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_237
timestamp 1704896540
transform 1 0 22908 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_245
timestamp 1704896540
transform 1 0 23644 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1704896540
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1704896540
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 1704896540
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_29
timestamp 1704896540
transform 1 0 3772 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_37
timestamp 1704896540
transform 1 0 4508 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_65
timestamp 1704896540
transform 1 0 7084 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_72
timestamp 1704896540
transform 1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_85
timestamp 1704896540
transform 1 0 8924 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_98
timestamp 1704896540
transform 1 0 10120 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_108
timestamp 1704896540
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_127
timestamp 1704896540
transform 1 0 12788 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_135
timestamp 1704896540
transform 1 0 13524 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1704896540
transform 1 0 13892 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_149
timestamp 1704896540
transform 1 0 14812 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_156
timestamp 1704896540
transform 1 0 15456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_163
timestamp 1704896540
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1704896540
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_175
timestamp 1704896540
transform 1 0 17204 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_183
timestamp 1704896540
transform 1 0 17940 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_205
timestamp 1704896540
transform 1 0 19964 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_215
timestamp 1704896540
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1704896540
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1704896540
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_237
timestamp 1704896540
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_245
timestamp 1704896540
transform 1 0 23644 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform -1 0 5796 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 11408 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 7268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 21620 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 4692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 3680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 7912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform -1 0 14812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform -1 0 16468 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 23368 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 21528 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform -1 0 23276 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform -1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform -1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 20240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform -1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 6164 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 18492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform -1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 12236 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 23736 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform -1 0 11408 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform -1 0 10120 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform -1 0 18584 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform 1 0 15088 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform 1 0 7544 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform 1 0 15640 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform -1 0 3680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform -1 0 9844 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform -1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform -1 0 19136 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform -1 0 18492 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform -1 0 10120 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 17112 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform -1 0 17848 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform -1 0 7084 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform -1 0 3956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 21712 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform -1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform -1 0 15548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform -1 0 21436 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 19964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform -1 0 6440 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform -1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform -1 0 8004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform 1 0 3864 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform -1 0 20240 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform 1 0 18584 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 21252 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform -1 0 10120 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform -1 0 18768 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform -1 0 23644 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform -1 0 11408 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform -1 0 15456 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform -1 0 14536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 16008 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform -1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform -1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform -1 0 13064 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1704896540
transform -1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform -1 0 23460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform -1 0 20240 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform -1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1704896540
transform -1 0 21896 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform -1 0 16376 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform -1 0 12236 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform -1 0 16836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform 1 0 19504 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1704896540
transform -1 0 21252 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform 1 0 20056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1704896540
transform -1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform -1 0 7912 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1704896540
transform 1 0 14168 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1704896540
transform -1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform -1 0 7084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform -1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1704896540
transform -1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1704896540
transform 1 0 23000 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform -1 0 12512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1704896540
transform -1 0 12236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform -1 0 18768 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1704896540
transform -1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform -1 0 12236 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform -1 0 16560 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform -1 0 6256 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform 1 0 8372 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform -1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform -1 0 21620 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform -1 0 18216 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform -1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1704896540
transform -1 0 6256 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1704896540
transform -1 0 22540 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1704896540
transform -1 0 18676 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1704896540
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1704896540
transform -1 0 5704 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1704896540
transform -1 0 11500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1704896540
transform -1 0 18216 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1704896540
transform -1 0 21436 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1704896540
transform -1 0 7544 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1704896540
transform -1 0 19964 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1704896540
transform -1 0 16836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1704896540
transform -1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1704896540
transform -1 0 20424 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1704896540
transform -1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1704896540
transform -1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1704896540
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1704896540
transform -1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1704896540
transform -1 0 18860 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1704896540
transform -1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1704896540
transform -1 0 22908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1704896540
transform -1 0 12696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform 1 0 8004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 9108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 12972 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 13616 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 20608 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1704896540
transform -1 0 23736 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1704896540
transform -1 0 20976 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1704896540
transform -1 0 23736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1704896540
transform -1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform -1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1704896540
transform -1 0 23736 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1704896540
transform -1 0 23736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1704896540
transform -1 0 23460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1704896540
transform 1 0 16192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1704896540
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1704896540
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1704896540
transform -1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1704896540
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1704896540
transform 1 0 13248 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1704896540
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1704896540
transform -1 0 5612 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1704896540
transform -1 0 4968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1704896540
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1704896540
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1704896540
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1704896540
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1704896540
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1704896540
transform -1 0 8832 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1704896540
transform 1 0 12236 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1704896540
transform -1 0 15456 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1704896540
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1704896540
transform -1 0 20608 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1704896540
transform -1 0 16100 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1704896540
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1704896540
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1704896540
transform 1 0 23368 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1704896540
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1704896540
transform -1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1704896540
transform 1 0 23368 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1704896540
transform 1 0 23368 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1704896540
transform 1 0 23368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1704896540
transform 1 0 23368 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1704896540
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 1704896540
transform -1 0 18032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1704896540
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output56
timestamp 1704896540
transform -1 0 17388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1704896540
transform 1 0 23368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1704896540
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1704896540
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1704896540
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1704896540
transform -1 0 12880 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1704896540
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1704896540
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1704896540
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output65
timestamp 1704896540
transform -1 0 11960 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1704896540
transform -1 0 6256 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1704896540
transform 1 0 7176 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1704896540
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1704896540
transform -1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1704896540
transform 1 0 6532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1704896540
transform -1 0 8832 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1704896540
transform -1 0 10580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1704896540
transform -1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 24012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 24012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 24012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 24012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 1704896540
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 24012 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 1704896540
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 1704896540
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 24012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 1704896540
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 1704896540
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 1704896540
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 1704896540
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 24012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 1704896540
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1704896540
transform -1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 1704896540
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1704896540
transform -1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 1704896540
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1704896540
transform -1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 1704896540
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1704896540
transform -1 0 24012 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 1704896540
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1704896540
transform -1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 1704896540
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1704896540
transform -1 0 24012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1704896540
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 1704896540
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 1704896540
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1704896540
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1704896540
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1704896540
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1704896540
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 1704896540
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 1704896540
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 1704896540
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 1704896540
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1704896540
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1704896540
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 1704896540
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1704896540
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1704896540
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1704896540
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1704896540
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1704896540
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 1704896540
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 1704896540
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 1704896540
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 1704896540
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1704896540
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1704896540
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 1704896540
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 1704896540
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1704896540
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1704896540
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 1704896540
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 1704896540
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1704896540
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1704896540
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 1704896540
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 1704896540
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1704896540
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1704896540
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 1704896540
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 1704896540
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1704896540
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1704896540
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 1704896540
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1704896540
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1704896540
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1704896540
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1704896540
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1704896540
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1704896540
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1704896540
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 1704896540
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 1704896540
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1704896540
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1704896540
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 1704896540
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 1704896540
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1704896540
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1704896540
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 1704896540
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 1704896540
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1704896540
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1704896540
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 1704896540
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 1704896540
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1704896540
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1704896540
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 1704896540
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 1704896540
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1704896540
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1704896540
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1704896540
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1704896540
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 1704896540
transform 1 0 3680 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 1704896540
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 1704896540
transform 1 0 8832 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 1704896540
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 1704896540
transform 1 0 13984 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 1704896540
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 1704896540
transform 1 0 19136 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 1704896540
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 23128 400 23248 0 FreeSans 480 0 0 0 Clk
port 0 nsew signal input
flabel metal3 s 0 13608 400 13728 0 FreeSans 480 0 0 0 Data_In[0]
port 1 nsew signal input
flabel metal2 s 8390 26924 8446 27324 0 FreeSans 224 90 0 0 Data_In[10]
port 2 nsew signal input
flabel metal2 s 9678 26924 9734 27324 0 FreeSans 224 90 0 0 Data_In[11]
port 3 nsew signal input
flabel metal2 s 12898 26924 12954 27324 0 FreeSans 224 90 0 0 Data_In[12]
port 4 nsew signal input
flabel metal2 s 14186 26924 14242 27324 0 FreeSans 224 90 0 0 Data_In[13]
port 5 nsew signal input
flabel metal2 s 18694 26924 18750 27324 0 FreeSans 224 90 0 0 Data_In[14]
port 6 nsew signal input
flabel metal2 s 13542 26924 13598 27324 0 FreeSans 224 90 0 0 Data_In[15]
port 7 nsew signal input
flabel metal2 s 19338 26924 19394 27324 0 FreeSans 224 90 0 0 Data_In[16]
port 8 nsew signal input
flabel metal3 s 24780 19728 25180 19848 0 FreeSans 480 0 0 0 Data_In[17]
port 9 nsew signal input
flabel metal3 s 24780 11568 25180 11688 0 FreeSans 480 0 0 0 Data_In[18]
port 10 nsew signal input
flabel metal3 s 24780 13608 25180 13728 0 FreeSans 480 0 0 0 Data_In[19]
port 11 nsew signal input
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 Data_In[1]
port 12 nsew signal input
flabel metal3 s 24780 14968 25180 15088 0 FreeSans 480 0 0 0 Data_In[20]
port 13 nsew signal input
flabel metal3 s 24780 17688 25180 17808 0 FreeSans 480 0 0 0 Data_In[21]
port 14 nsew signal input
flabel metal3 s 24780 17008 25180 17128 0 FreeSans 480 0 0 0 Data_In[22]
port 15 nsew signal input
flabel metal3 s 24780 10888 25180 11008 0 FreeSans 480 0 0 0 Data_In[23]
port 16 nsew signal input
flabel metal3 s 24780 8848 25180 8968 0 FreeSans 480 0 0 0 Data_In[24]
port 17 nsew signal input
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 Data_In[25]
port 18 nsew signal input
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 Data_In[26]
port 19 nsew signal input
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 Data_In[27]
port 20 nsew signal input
flabel metal3 s 24780 6128 25180 6248 0 FreeSans 480 0 0 0 Data_In[28]
port 21 nsew signal input
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 Data_In[29]
port 22 nsew signal input
flabel metal3 s 0 8848 400 8968 0 FreeSans 480 0 0 0 Data_In[2]
port 23 nsew signal input
flabel metal2 s 12254 26924 12310 27324 0 FreeSans 224 90 0 0 Data_In[30]
port 24 nsew signal input
flabel metal3 s 0 12248 400 12368 0 FreeSans 480 0 0 0 Data_In[31]
port 25 nsew signal input
flabel metal3 s 0 11568 400 11688 0 FreeSans 480 0 0 0 Data_In[3]
port 26 nsew signal input
flabel metal3 s 0 14968 400 15088 0 FreeSans 480 0 0 0 Data_In[4]
port 27 nsew signal input
flabel metal3 s 0 15648 400 15768 0 FreeSans 480 0 0 0 Data_In[5]
port 28 nsew signal input
flabel metal2 s 9034 26924 9090 27324 0 FreeSans 224 90 0 0 Data_In[6]
port 29 nsew signal input
flabel metal2 s 5814 26924 5870 27324 0 FreeSans 224 90 0 0 Data_In[7]
port 30 nsew signal input
flabel metal2 s 5170 26924 5226 27324 0 FreeSans 224 90 0 0 Data_In[8]
port 31 nsew signal input
flabel metal3 s 0 18368 400 18488 0 FreeSans 480 0 0 0 Data_In[9]
port 32 nsew signal input
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 FClrN
port 33 nsew signal input
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 FInN
port 34 nsew signal input
flabel metal2 s 9034 0 9090 400 0 FreeSans 224 90 0 0 FOutN
port 35 nsew signal input
flabel metal3 s 0 12928 400 13048 0 FreeSans 480 0 0 0 F_Data[0]
port 36 nsew signal output
flabel metal2 s 10322 26924 10378 27324 0 FreeSans 224 90 0 0 F_Data[10]
port 37 nsew signal output
flabel metal2 s 11610 26924 11666 27324 0 FreeSans 224 90 0 0 F_Data[11]
port 38 nsew signal output
flabel metal2 s 14830 26924 14886 27324 0 FreeSans 224 90 0 0 F_Data[12]
port 39 nsew signal output
flabel metal2 s 16118 26924 16174 27324 0 FreeSans 224 90 0 0 F_Data[13]
port 40 nsew signal output
flabel metal2 s 19982 26924 20038 27324 0 FreeSans 224 90 0 0 F_Data[14]
port 41 nsew signal output
flabel metal2 s 15474 26924 15530 27324 0 FreeSans 224 90 0 0 F_Data[15]
port 42 nsew signal output
flabel metal3 s 24780 21088 25180 21208 0 FreeSans 480 0 0 0 F_Data[16]
port 43 nsew signal output
flabel metal3 s 24780 18368 25180 18488 0 FreeSans 480 0 0 0 F_Data[17]
port 44 nsew signal output
flabel metal3 s 24780 12248 25180 12368 0 FreeSans 480 0 0 0 F_Data[18]
port 45 nsew signal output
flabel metal3 s 24780 12928 25180 13048 0 FreeSans 480 0 0 0 F_Data[19]
port 46 nsew signal output
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 F_Data[1]
port 47 nsew signal output
flabel metal3 s 24780 16328 25180 16448 0 FreeSans 480 0 0 0 F_Data[20]
port 48 nsew signal output
flabel metal3 s 24780 19048 25180 19168 0 FreeSans 480 0 0 0 F_Data[21]
port 49 nsew signal output
flabel metal3 s 24780 15648 25180 15768 0 FreeSans 480 0 0 0 F_Data[22]
port 50 nsew signal output
flabel metal3 s 24780 10208 25180 10328 0 FreeSans 480 0 0 0 F_Data[23]
port 51 nsew signal output
flabel metal3 s 24780 9528 25180 9648 0 FreeSans 480 0 0 0 F_Data[24]
port 52 nsew signal output
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 F_Data[25]
port 53 nsew signal output
flabel metal2 s 21270 0 21326 400 0 FreeSans 224 90 0 0 F_Data[26]
port 54 nsew signal output
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 F_Data[27]
port 55 nsew signal output
flabel metal3 s 24780 6808 25180 6928 0 FreeSans 480 0 0 0 F_Data[28]
port 56 nsew signal output
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 F_Data[29]
port 57 nsew signal output
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 F_Data[2]
port 58 nsew signal output
flabel metal3 s 24780 14288 25180 14408 0 FreeSans 480 0 0 0 F_Data[30]
port 59 nsew signal output
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 F_Data[31]
port 60 nsew signal output
flabel metal3 s 0 10888 400 11008 0 FreeSans 480 0 0 0 F_Data[3]
port 61 nsew signal output
flabel metal3 s 0 14288 400 14408 0 FreeSans 480 0 0 0 F_Data[4]
port 62 nsew signal output
flabel metal3 s 0 16328 400 16448 0 FreeSans 480 0 0 0 F_Data[5]
port 63 nsew signal output
flabel metal2 s 10966 26924 11022 27324 0 FreeSans 224 90 0 0 F_Data[6]
port 64 nsew signal output
flabel metal2 s 6458 26924 6514 27324 0 FreeSans 224 90 0 0 F_Data[7]
port 65 nsew signal output
flabel metal2 s 7102 26924 7158 27324 0 FreeSans 224 90 0 0 F_Data[8]
port 66 nsew signal output
flabel metal3 s 0 19048 400 19168 0 FreeSans 480 0 0 0 F_Data[9]
port 67 nsew signal output
flabel metal2 s 7102 0 7158 400 0 FreeSans 224 90 0 0 F_EmptyN
port 68 nsew signal output
flabel metal2 s 6458 0 6514 400 0 FreeSans 224 90 0 0 F_FirstN
port 69 nsew signal output
flabel metal2 s 8390 0 8446 400 0 FreeSans 224 90 0 0 F_FullN
port 70 nsew signal output
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 F_LastN
port 71 nsew signal output
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 F_SLastN
port 72 nsew signal output
flabel metal2 s 5814 0 5870 400 0 FreeSans 224 90 0 0 RstN
port 73 nsew signal input
flabel metal4 s 2844 2128 3164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 5844 2128 6164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 8844 2128 9164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 11844 2128 12164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 14844 2128 15164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 17844 2128 18164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 20844 2128 21164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 23844 2128 24164 25072 0 FreeSans 1920 90 0 0 VGND
port 74 nsew ground bidirectional
flabel metal4 s 1344 2128 1664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 4344 2128 4664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 7344 2128 7664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 10344 2128 10664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 13344 2128 13664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 16344 2128 16664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 19344 2128 19664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
flabel metal4 s 22344 2128 22664 25072 0 FreeSans 1920 90 0 0 VPWR
port 75 nsew power bidirectional
rlabel metal1 12634 25024 12634 25024 0 VGND
rlabel metal1 12558 24480 12558 24480 0 VPWR
rlabel metal3 1855 23188 1855 23188 0 Clk
rlabel metal3 774 13668 774 13668 0 Data_In[0]
rlabel metal1 8234 24786 8234 24786 0 Data_In[10]
rlabel metal1 9430 24786 9430 24786 0 Data_In[11]
rlabel metal1 12972 24786 12972 24786 0 Data_In[12]
rlabel metal1 14398 24174 14398 24174 0 Data_In[13]
rlabel metal1 18860 24786 18860 24786 0 Data_In[14]
rlabel metal1 13616 24786 13616 24786 0 Data_In[15]
rlabel metal1 20654 24752 20654 24752 0 Data_In[16]
rlabel metal2 23690 20111 23690 20111 0 Data_In[17]
rlabel metal2 23506 11713 23506 11713 0 Data_In[18]
rlabel metal3 24296 13668 24296 13668 0 Data_In[19]
rlabel metal3 360 9588 360 9588 0 Data_In[1]
rlabel metal2 21574 14161 21574 14161 0 Data_In[20]
rlabel metal2 23322 19091 23322 19091 0 Data_In[21]
rlabel metal1 23736 19822 23736 19822 0 Data_In[22]
rlabel metal1 23690 8976 23690 8976 0 Data_In[23]
rlabel via2 23414 8925 23414 8925 0 Data_In[24]
rlabel metal2 16146 1384 16146 1384 0 Data_In[25]
rlabel metal2 19366 1384 19366 1384 0 Data_In[26]
rlabel metal2 15502 1384 15502 1384 0 Data_In[27]
rlabel metal2 23690 6239 23690 6239 0 Data_In[28]
rlabel metal2 14214 1384 14214 1384 0 Data_In[29]
rlabel metal3 360 8908 360 8908 0 Data_In[2]
rlabel metal2 12282 25850 12282 25850 0 Data_In[30]
rlabel metal3 360 12308 360 12308 0 Data_In[31]
rlabel metal3 360 11628 360 11628 0 Data_In[3]
rlabel metal3 866 15028 866 15028 0 Data_In[4]
rlabel metal3 544 15708 544 15708 0 Data_In[5]
rlabel metal1 8694 24174 8694 24174 0 Data_In[6]
rlabel metal2 5566 25585 5566 25585 0 Data_In[7]
rlabel metal1 5060 24786 5060 24786 0 Data_In[8]
rlabel metal3 360 18428 360 18428 0 Data_In[9]
rlabel metal2 10350 1384 10350 1384 0 FClrN
rlabel metal2 11638 1384 11638 1384 0 FInN
rlabel metal2 9062 823 9062 823 0 FOutN
rlabel metal1 1426 12954 1426 12954 0 F_Data[0]
rlabel metal1 9430 24650 9430 24650 0 F_Data[10]
rlabel metal2 11638 25782 11638 25782 0 F_Data[11]
rlabel metal1 14858 24786 14858 24786 0 F_Data[12]
rlabel metal1 16514 24582 16514 24582 0 F_Data[13]
rlabel metal1 20056 24786 20056 24786 0 F_Data[14]
rlabel metal1 15548 24786 15548 24786 0 F_Data[15]
rlabel metal3 24250 21148 24250 21148 0 F_Data[16]
rlabel metal3 24618 18428 24618 18428 0 F_Data[17]
rlabel via2 23598 12325 23598 12325 0 F_Data[18]
rlabel metal3 24618 12988 24618 12988 0 F_Data[19]
rlabel metal3 659 10268 659 10268 0 F_Data[1]
rlabel metal3 24641 16388 24641 16388 0 F_Data[20]
rlabel metal3 24250 19108 24250 19108 0 F_Data[21]
rlabel metal1 23506 15130 23506 15130 0 F_Data[22]
rlabel metal1 23506 9418 23506 9418 0 F_Data[23]
rlabel metal3 23882 9588 23882 9588 0 F_Data[24]
rlabel metal2 17434 1350 17434 1350 0 F_Data[25]
rlabel metal2 21298 1316 21298 1316 0 F_Data[26]
rlabel metal2 16790 1350 16790 1350 0 F_Data[27]
rlabel metal3 24158 6868 24158 6868 0 F_Data[28]
rlabel metal2 14858 755 14858 755 0 F_Data[29]
rlabel metal3 774 8228 774 8228 0 F_Data[2]
rlabel metal3 24250 14348 24250 14348 0 F_Data[30]
rlabel metal2 12282 1350 12282 1350 0 F_Data[31]
rlabel metal3 912 10948 912 10948 0 F_Data[3]
rlabel metal3 544 14348 544 14348 0 F_Data[4]
rlabel metal1 1426 16422 1426 16422 0 F_Data[5]
rlabel metal1 11270 24378 11270 24378 0 F_Data[6]
rlabel metal1 6256 24582 6256 24582 0 F_Data[7]
rlabel metal1 7268 24582 7268 24582 0 F_Data[8]
rlabel metal3 774 19108 774 19108 0 F_Data[9]
rlabel metal2 7130 1350 7130 1350 0 F_EmptyN
rlabel metal2 6486 1316 6486 1316 0 F_FirstN
rlabel metal2 8418 1316 8418 1316 0 F_FullN
rlabel metal2 9706 1350 9706 1350 0 F_LastN
rlabel metal2 7774 1350 7774 1350 0 F_SLastN
rlabel metal2 5842 823 5842 823 0 RstN
rlabel metal2 1886 13090 1886 13090 0 _000_
rlabel metal2 6486 10098 6486 10098 0 _001_
rlabel metal2 3358 8024 3358 8024 0 _002_
rlabel metal1 1886 9690 1886 9690 0 _003_
rlabel metal1 6568 12818 6568 12818 0 _004_
rlabel metal2 2898 15912 2898 15912 0 _005_
rlabel metal1 8413 20502 8413 20502 0 _006_
rlabel metal2 3450 23970 3450 23970 0 _007_
rlabel via1 3537 20434 3537 20434 0 _008_
rlabel metal1 3629 18326 3629 18326 0 _009_
rlabel metal1 7861 16558 7861 16558 0 _010_
rlabel metal2 8326 23528 8326 23528 0 _011_
rlabel metal2 12558 18462 12558 18462 0 _012_
rlabel metal1 12512 21862 12512 21862 0 _013_
rlabel metal2 17158 22882 17158 22882 0 _014_
rlabel metal2 12558 23562 12558 23562 0 _015_
rlabel metal1 16744 20298 16744 20298 0 _016_
rlabel metal1 16785 17578 16785 17578 0 _017_
rlabel metal1 14664 12206 14664 12206 0 _018_
rlabel metal1 19458 12614 19458 12614 0 _019_
rlabel metal2 20010 14790 20010 14790 0 _020_
rlabel metal1 20332 17306 20332 17306 0 _021_
rlabel metal2 15226 14178 15226 14178 0 _022_
rlabel metal1 19780 10234 19780 10234 0 _023_
rlabel metal2 16330 8738 16330 8738 0 _024_
rlabel metal1 14204 5678 14204 5678 0 _025_
rlabel metal1 18262 2618 18262 2618 0 _026_
rlabel metal1 14398 3706 14398 3706 0 _027_
rlabel metal2 18998 6086 18998 6086 0 _028_
rlabel metal1 12732 8942 12732 8942 0 _029_
rlabel metal1 10212 14586 10212 14586 0 _030_
rlabel via1 9425 11730 9425 11730 0 _031_
rlabel metal1 11684 6358 11684 6358 0 _032_
rlabel metal1 10304 7922 10304 7922 0 _033_
rlabel metal2 4416 12716 4416 12716 0 _034_
rlabel metal1 7482 9962 7482 9962 0 _035_
rlabel metal1 4446 7786 4446 7786 0 _036_
rlabel via1 4926 9962 4926 9962 0 _037_
rlabel metal1 9614 14586 9614 14586 0 _038_
rlabel via1 5101 15470 5101 15470 0 _039_
rlabel metal1 9890 20536 9890 20536 0 _040_
rlabel metal1 7410 23766 7410 23766 0 _041_
rlabel metal1 8004 21862 8004 21862 0 _042_
rlabel metal1 7544 17850 7544 17850 0 _043_
rlabel metal1 9690 18326 9690 18326 0 _044_
rlabel metal1 9920 23766 9920 23766 0 _045_
rlabel via1 14853 17578 14853 17578 0 _046_
rlabel metal2 16146 20774 16146 20774 0 _047_
rlabel metal1 19688 22746 19688 22746 0 _048_
rlabel metal1 16652 23834 16652 23834 0 _049_
rlabel metal1 20056 20570 20056 20570 0 _050_
rlabel metal1 20336 17578 20336 17578 0 _051_
rlabel via1 17429 11798 17429 11798 0 _052_
rlabel metal1 21988 12410 21988 12410 0 _053_
rlabel metal2 21482 14824 21482 14824 0 _054_
rlabel metal1 22857 17238 22857 17238 0 _055_
rlabel metal1 17424 14382 17424 14382 0 _056_
rlabel metal2 22126 9996 22126 9996 0 _057_
rlabel metal1 19504 8602 19504 8602 0 _058_
rlabel metal2 16238 5984 16238 5984 0 _059_
rlabel metal2 21298 4386 21298 4386 0 _060_
rlabel metal1 17204 3978 17204 3978 0 _061_
rlabel metal1 21932 6766 21932 6766 0 _062_
rlabel metal1 14950 8602 14950 8602 0 _063_
rlabel via1 12829 14382 12829 14382 0 _064_
rlabel metal2 11362 13022 11362 13022 0 _065_
rlabel via1 3537 13906 3537 13906 0 _066_
rlabel metal1 6992 10778 6992 10778 0 _067_
rlabel metal1 4124 7446 4124 7446 0 _068_
rlabel metal1 3848 11050 3848 11050 0 _069_
rlabel metal1 7824 14382 7824 14382 0 _070_
rlabel metal2 5290 15640 5290 15640 0 _071_
rlabel metal1 10299 20502 10299 20502 0 _072_
rlabel metal1 5428 23834 5428 23834 0 _073_
rlabel metal1 5474 22406 5474 22406 0 _074_
rlabel via1 5653 17578 5653 17578 0 _075_
rlabel metal2 10258 16966 10258 16966 0 _076_
rlabel metal2 9890 23970 9890 23970 0 _077_
rlabel via1 13565 17238 13565 17238 0 _078_
rlabel metal1 14112 20434 14112 20434 0 _079_
rlabel metal1 19258 23018 19258 23018 0 _080_
rlabel via1 14393 23018 14393 23018 0 _081_
rlabel metal1 19596 20026 19596 20026 0 _082_
rlabel metal1 18487 17238 18487 17238 0 _083_
rlabel via1 17153 12206 17153 12206 0 _084_
rlabel via1 22121 12206 22121 12206 0 _085_
rlabel metal1 23184 14042 23184 14042 0 _086_
rlabel metal2 21850 18632 21850 18632 0 _087_
rlabel metal1 16866 15062 16866 15062 0 _088_
rlabel via1 21201 8942 21201 8942 0 _089_
rlabel metal1 17756 8058 17756 8058 0 _090_
rlabel metal1 16932 6358 16932 6358 0 _091_
rlabel metal1 21129 3434 21129 3434 0 _092_
rlabel metal1 15962 3128 15962 3128 0 _093_
rlabel metal2 21390 6902 21390 6902 0 _094_
rlabel metal1 13064 11322 13064 11322 0 _095_
rlabel metal2 12466 15266 12466 15266 0 _096_
rlabel via1 13202 13413 13202 13413 0 _097_
rlabel via1 1881 13906 1881 13906 0 _098_
rlabel via1 6766 10030 6766 10030 0 _099_
rlabel metal1 2203 8534 2203 8534 0 _100_
rlabel metal1 1973 10710 1973 10710 0 _101_
rlabel via1 6205 13294 6205 13294 0 _102_
rlabel metal1 2484 16218 2484 16218 0 _103_
rlabel metal1 8924 21114 8924 21114 0 _104_
rlabel metal1 3864 23290 3864 23290 0 _105_
rlabel metal2 3818 21318 3818 21318 0 _106_
rlabel metal1 3496 18938 3496 18938 0 _107_
rlabel metal2 7774 17442 7774 17442 0 _108_
rlabel metal1 8321 22678 8321 22678 0 _109_
rlabel metal1 12180 17646 12180 17646 0 _110_
rlabel metal2 12742 21182 12742 21182 0 _111_
rlabel metal2 16882 23426 16882 23426 0 _112_
rlabel metal1 12645 23766 12645 23766 0 _113_
rlabel metal1 16744 21114 16744 21114 0 _114_
rlabel metal1 16836 17306 16836 17306 0 _115_
rlabel viali 14853 12818 14853 12818 0 _116_
rlabel via1 19453 12818 19453 12818 0 _117_
rlabel metal1 19729 15402 19729 15402 0 _118_
rlabel via1 20465 18734 20465 18734 0 _119_
rlabel via1 15129 15470 15129 15470 0 _120_
rlabel metal2 20102 10642 20102 10642 0 _121_
rlabel metal1 16606 9690 16606 9690 0 _122_
rlabel metal1 14296 6290 14296 6290 0 _123_
rlabel metal1 18395 3094 18395 3094 0 _124_
rlabel via1 13749 3026 13749 3026 0 _125_
rlabel metal2 18538 6086 18538 6086 0 _126_
rlabel metal1 13100 9554 13100 9554 0 _127_
rlabel metal1 11219 14314 11219 14314 0 _128_
rlabel metal1 9476 12614 9476 12614 0 _129_
rlabel metal2 6854 7565 6854 7565 0 _130_
rlabel metal1 9936 5882 9936 5882 0 _131_
rlabel metal1 6716 6834 6716 6834 0 _132_
rlabel metal1 5750 5338 5750 5338 0 _133_
rlabel metal2 5566 3740 5566 3740 0 _134_
rlabel metal1 6946 3128 6946 3128 0 _135_
rlabel metal1 12052 2618 12052 2618 0 _136_
rlabel metal2 13202 3298 13202 3298 0 _137_
rlabel metal2 10810 9180 10810 9180 0 _138_
rlabel metal2 10534 9826 10534 9826 0 _139_
rlabel metal2 13294 15436 13294 15436 0 _140_
rlabel metal1 4416 13362 4416 13362 0 _141_
rlabel metal2 12742 15742 12742 15742 0 _142_
rlabel metal1 5520 13362 5520 13362 0 _143_
rlabel metal1 5704 13498 5704 13498 0 _144_
rlabel metal1 7682 10438 7682 10438 0 _145_
rlabel metal1 5842 8534 5842 8534 0 _146_
rlabel metal1 5336 10778 5336 10778 0 _147_
rlabel metal1 9384 13906 9384 13906 0 _148_
rlabel metal2 6624 23052 6624 23052 0 _149_
rlabel metal2 5658 22100 5658 22100 0 _150_
rlabel metal1 6762 16660 6762 16660 0 _151_
rlabel metal2 11178 20332 11178 20332 0 _152_
rlabel metal1 8050 23188 8050 23188 0 _153_
rlabel metal1 6946 19822 6946 19822 0 _154_
rlabel metal1 5428 18938 5428 18938 0 _155_
rlabel metal1 10120 17850 10120 17850 0 _156_
rlabel metal1 14904 18122 14904 18122 0 _157_
rlabel metal1 14720 18190 14720 18190 0 _158_
rlabel metal1 11132 23290 11132 23290 0 _159_
rlabel metal1 13800 18190 13800 18190 0 _160_
rlabel metal1 16008 20910 16008 20910 0 _161_
rlabel metal1 21666 23732 21666 23732 0 _162_
rlabel metal2 13938 23936 13938 23936 0 _163_
rlabel metal1 20378 20332 20378 20332 0 _164_
rlabel metal1 18538 15606 18538 15606 0 _165_
rlabel metal2 22034 16915 22034 16915 0 _166_
rlabel metal1 19734 18258 19734 18258 0 _167_
rlabel metal1 18630 12886 18630 12886 0 _168_
rlabel metal1 21896 12614 21896 12614 0 _169_
rlabel metal1 21206 15674 21206 15674 0 _170_
rlabel metal2 22586 18445 22586 18445 0 _171_
rlabel metal1 18538 15402 18538 15402 0 _172_
rlabel metal1 18952 9418 18952 9418 0 _173_
rlabel metal1 20102 4046 20102 4046 0 _174_
rlabel metal1 22724 8942 22724 8942 0 _175_
rlabel metal1 20654 9588 20654 9588 0 _176_
rlabel metal1 16698 5542 16698 5542 0 _177_
rlabel metal1 22126 3536 22126 3536 0 _178_
rlabel metal1 17434 3026 17434 3026 0 _179_
rlabel metal1 21574 6290 21574 6290 0 _180_
rlabel metal2 14122 10438 14122 10438 0 _181_
rlabel metal2 14306 14620 14306 14620 0 _182_
rlabel metal1 12328 12818 12328 12818 0 _183_
rlabel metal2 12650 8143 12650 8143 0 _184_
rlabel metal2 14214 16677 14214 16677 0 _185_
rlabel metal1 6302 12614 6302 12614 0 _186_
rlabel metal1 2116 12818 2116 12818 0 _187_
rlabel metal2 6670 9146 6670 9146 0 _188_
rlabel metal1 3450 7514 3450 7514 0 _189_
rlabel metal1 2300 9554 2300 9554 0 _190_
rlabel metal1 6026 12886 6026 12886 0 _191_
rlabel metal1 3312 15470 3312 15470 0 _192_
rlabel metal2 4922 22372 4922 22372 0 _193_
rlabel metal1 8878 20026 8878 20026 0 _194_
rlabel metal2 4278 23256 4278 23256 0 _195_
rlabel metal2 4738 21488 4738 21488 0 _196_
rlabel metal1 4094 18734 4094 18734 0 _197_
rlabel metal1 8372 17170 8372 17170 0 _198_
rlabel metal1 8740 23086 8740 23086 0 _199_
rlabel metal1 17664 19890 17664 19890 0 _200_
rlabel metal1 12880 18734 12880 18734 0 _201_
rlabel metal2 14030 21794 14030 21794 0 _202_
rlabel metal2 17342 23052 17342 23052 0 _203_
rlabel metal1 12006 24140 12006 24140 0 _204_
rlabel metal2 17250 20196 17250 20196 0 _205_
rlabel metal1 17756 17850 17756 17850 0 _206_
rlabel metal1 16192 16014 16192 16014 0 _207_
rlabel metal1 15916 12886 15916 12886 0 _208_
rlabel metal1 18998 12818 18998 12818 0 _209_
rlabel metal1 20516 14382 20516 14382 0 _210_
rlabel metal1 20516 17170 20516 17170 0 _211_
rlabel metal2 15410 14892 15410 14892 0 _212_
rlabel metal1 20010 10064 20010 10064 0 _213_
rlabel metal1 15594 2924 15594 2924 0 _214_
rlabel metal1 16514 8500 16514 8500 0 _215_
rlabel metal2 13846 6460 13846 6460 0 _216_
rlabel metal1 18814 2414 18814 2414 0 _217_
rlabel metal1 15088 3162 15088 3162 0 _218_
rlabel metal2 18814 6426 18814 6426 0 _219_
rlabel metal2 12558 9724 12558 9724 0 _220_
rlabel metal1 10396 14382 10396 14382 0 _221_
rlabel metal1 9338 11322 9338 11322 0 _222_
rlabel metal1 11868 6698 11868 6698 0 _223_
rlabel metal2 12742 7616 12742 7616 0 _224_
rlabel metal1 12512 5610 12512 5610 0 _225_
rlabel metal1 12328 5882 12328 5882 0 _226_
rlabel metal1 11500 6766 11500 6766 0 _227_
rlabel metal2 15686 10234 15686 10234 0 _228_
rlabel metal1 13524 13362 13524 13362 0 _229_
rlabel metal1 4692 14450 4692 14450 0 _230_
rlabel metal1 11914 7514 11914 7514 0 _231_
rlabel via1 7958 7837 7958 7837 0 _232_
rlabel metal1 14398 7854 14398 7854 0 _233_
rlabel metal1 16606 16082 16606 16082 0 _234_
rlabel metal1 6808 16014 6808 16014 0 _235_
rlabel metal1 4094 13974 4094 13974 0 _236_
rlabel metal1 7268 9690 7268 9690 0 _237_
rlabel metal1 4140 7854 4140 7854 0 _238_
rlabel metal1 3772 9690 3772 9690 0 _239_
rlabel metal1 9982 14348 9982 14348 0 _240_
rlabel metal1 5980 15878 5980 15878 0 _241_
rlabel metal1 6302 23528 6302 23528 0 _242_
rlabel metal1 9936 20026 9936 20026 0 _243_
rlabel metal2 7130 24004 7130 24004 0 _244_
rlabel metal1 7452 20570 7452 20570 0 _245_
rlabel metal2 7130 17850 7130 17850 0 _246_
rlabel metal2 9338 18428 9338 18428 0 _247_
rlabel metal1 9476 23698 9476 23698 0 _248_
rlabel metal1 19826 18870 19826 18870 0 _249_
rlabel metal1 15502 18394 15502 18394 0 _250_
rlabel metal2 15962 20026 15962 20026 0 _251_
rlabel metal2 18906 23324 18906 23324 0 _252_
rlabel metal1 16560 23290 16560 23290 0 _253_
rlabel metal1 20286 20468 20286 20468 0 _254_
rlabel metal1 18998 18734 18998 18734 0 _255_
rlabel metal2 18998 15402 18998 15402 0 _256_
rlabel metal1 17572 13294 17572 13294 0 _257_
rlabel metal1 21712 13158 21712 13158 0 _258_
rlabel metal2 20838 15674 20838 15674 0 _259_
rlabel metal1 22954 16422 22954 16422 0 _260_
rlabel metal1 17572 14994 17572 14994 0 _261_
rlabel metal2 21482 10404 21482 10404 0 _262_
rlabel metal1 17388 2958 17388 2958 0 _263_
rlabel metal2 19274 8262 19274 8262 0 _264_
rlabel metal1 16284 5202 16284 5202 0 _265_
rlabel metal1 21160 3162 21160 3162 0 _266_
rlabel metal2 17434 3638 17434 3638 0 _267_
rlabel metal1 21068 5882 21068 5882 0 _268_
rlabel metal2 15318 8908 15318 8908 0 _269_
rlabel metal2 14030 15606 14030 15606 0 _270_
rlabel metal1 11362 11866 11362 11866 0 _271_
rlabel metal1 3726 14382 3726 14382 0 _272_
rlabel metal1 6946 10642 6946 10642 0 _273_
rlabel metal2 3818 7956 3818 7956 0 _274_
rlabel metal2 3450 11322 3450 11322 0 _275_
rlabel metal1 7176 14994 7176 14994 0 _276_
rlabel metal1 6900 22542 6900 22542 0 _277_
rlabel metal2 5474 15980 5474 15980 0 _278_
rlabel metal2 11546 21828 11546 21828 0 _279_
rlabel metal1 6348 22746 6348 22746 0 _280_
rlabel metal1 6210 22610 6210 22610 0 _281_
rlabel metal1 6118 18258 6118 18258 0 _282_
rlabel metal1 10672 16558 10672 16558 0 _283_
rlabel metal1 11178 22474 11178 22474 0 _284_
rlabel metal1 10120 22746 10120 22746 0 _285_
rlabel metal2 14122 17204 14122 17204 0 _286_
rlabel metal1 14168 20026 14168 20026 0 _287_
rlabel metal1 18860 23086 18860 23086 0 _288_
rlabel metal1 14260 22746 14260 22746 0 _289_
rlabel metal1 19228 19822 19228 19822 0 _290_
rlabel metal1 22678 11662 22678 11662 0 _291_
rlabel metal1 18906 16762 18906 16762 0 _292_
rlabel metal1 17894 13362 17894 13362 0 _293_
rlabel metal1 21666 11866 21666 11866 0 _294_
rlabel metal1 23092 13906 23092 13906 0 _295_
rlabel metal1 22724 18938 22724 18938 0 _296_
rlabel metal1 16514 15470 16514 15470 0 _297_
rlabel metal1 20332 7922 20332 7922 0 _298_
rlabel metal1 21344 9554 21344 9554 0 _299_
rlabel metal1 17756 7854 17756 7854 0 _300_
rlabel metal1 16744 5338 16744 5338 0 _301_
rlabel metal1 21804 3502 21804 3502 0 _302_
rlabel metal2 15778 3468 15778 3468 0 _303_
rlabel metal2 21206 7004 21206 7004 0 _304_
rlabel metal1 13202 11152 13202 11152 0 _305_
rlabel metal1 12558 13498 12558 13498 0 _306_
rlabel metal1 10764 11866 10764 11866 0 _307_
rlabel metal1 14076 7854 14076 7854 0 _308_
rlabel metal1 13340 11254 13340 11254 0 _309_
rlabel metal1 7590 13838 7590 13838 0 _310_
rlabel metal1 2300 14382 2300 14382 0 _311_
rlabel metal1 6302 9690 6302 9690 0 _312_
rlabel metal1 2576 8942 2576 8942 0 _313_
rlabel metal1 2392 11118 2392 11118 0 _314_
rlabel metal2 6578 14212 6578 14212 0 _315_
rlabel metal2 2254 15844 2254 15844 0 _316_
rlabel metal1 5152 23154 5152 23154 0 _317_
rlabel metal1 9108 21862 9108 21862 0 _318_
rlabel metal1 4232 23086 4232 23086 0 _319_
rlabel metal1 4094 20910 4094 20910 0 _320_
rlabel metal1 4140 18394 4140 18394 0 _321_
rlabel metal1 7958 17136 7958 17136 0 _322_
rlabel metal1 8510 24140 8510 24140 0 _323_
rlabel metal1 16744 17034 16744 17034 0 _324_
rlabel metal2 12742 18700 12742 18700 0 _325_
rlabel metal2 13202 21828 13202 21828 0 _326_
rlabel metal1 17158 22610 17158 22610 0 _327_
rlabel metal1 13064 24174 13064 24174 0 _328_
rlabel metal1 16422 20876 16422 20876 0 _329_
rlabel metal1 17112 17170 17112 17170 0 _330_
rlabel metal1 20654 15980 20654 15980 0 _331_
rlabel metal1 15272 13294 15272 13294 0 _332_
rlabel metal1 20608 12954 20608 12954 0 _333_
rlabel metal1 20056 16082 20056 16082 0 _334_
rlabel via1 20746 19333 20746 19333 0 _335_
rlabel metal2 15594 15334 15594 15334 0 _336_
rlabel metal1 20516 10030 20516 10030 0 _337_
rlabel metal1 16146 6256 16146 6256 0 _338_
rlabel metal2 16790 9078 16790 9078 0 _339_
rlabel metal1 13570 6358 13570 6358 0 _340_
rlabel metal2 18906 3978 18906 3978 0 _341_
rlabel metal1 14076 3502 14076 3502 0 _342_
rlabel metal1 18538 5678 18538 5678 0 _343_
rlabel metal1 12650 9588 12650 9588 0 _344_
rlabel metal1 11546 14994 11546 14994 0 _345_
rlabel metal1 9798 12818 9798 12818 0 _346_
rlabel metal1 8648 7922 8648 7922 0 _347_
rlabel metal1 10718 4794 10718 4794 0 _348_
rlabel metal1 8878 6834 8878 6834 0 _349_
rlabel metal1 9200 7378 9200 7378 0 _350_
rlabel metal1 8096 8058 8096 8058 0 _351_
rlabel metal1 9476 7378 9476 7378 0 _352_
rlabel metal1 9338 6970 9338 6970 0 _353_
rlabel metal1 7912 4522 7912 4522 0 _354_
rlabel metal1 9384 3978 9384 3978 0 _355_
rlabel metal2 9798 6290 9798 6290 0 _356_
rlabel metal1 10120 5678 10120 5678 0 _357_
rlabel metal1 7912 6970 7912 6970 0 _358_
rlabel metal2 8418 4352 8418 4352 0 _359_
rlabel metal1 8740 3978 8740 3978 0 _360_
rlabel metal1 8326 7514 8326 7514 0 _361_
rlabel metal1 6578 5100 6578 5100 0 _362_
rlabel metal1 6624 4590 6624 4590 0 _363_
rlabel metal1 6118 5168 6118 5168 0 _364_
rlabel metal1 7958 4658 7958 4658 0 _365_
rlabel metal2 7038 5372 7038 5372 0 _366_
rlabel metal1 6670 4998 6670 4998 0 _367_
rlabel metal2 5750 4284 5750 4284 0 _368_
rlabel metal1 7406 4250 7406 4250 0 _369_
rlabel metal2 7222 4862 7222 4862 0 _370_
rlabel metal1 8970 4794 8970 4794 0 _371_
rlabel metal1 7130 4692 7130 4692 0 _372_
rlabel metal1 7728 3502 7728 3502 0 _373_
rlabel metal1 10396 4250 10396 4250 0 _374_
rlabel metal1 10626 3570 10626 3570 0 _375_
rlabel metal2 9522 3774 9522 3774 0 _376_
rlabel metal1 9522 3502 9522 3502 0 _377_
rlabel metal1 9798 3570 9798 3570 0 _378_
rlabel metal2 10902 2890 10902 2890 0 _379_
rlabel metal2 10994 3196 10994 3196 0 _380_
rlabel metal1 10672 2822 10672 2822 0 _381_
rlabel metal1 10488 3026 10488 3026 0 _382_
rlabel metal2 10718 3570 10718 3570 0 _383_
rlabel metal1 11362 3026 11362 3026 0 _384_
rlabel metal1 9430 9044 9430 9044 0 _385_
rlabel metal1 9300 8602 9300 8602 0 _386_
rlabel metal1 9936 8602 9936 8602 0 _387_
rlabel metal2 9706 9316 9706 9316 0 _388_
rlabel metal1 13800 14042 13800 14042 0 clknet_0_Clk
rlabel metal2 1886 8126 1886 8126 0 clknet_4_0_0_Clk
rlabel metal2 17802 3536 17802 3536 0 clknet_4_10_0_Clk
rlabel metal1 22218 10540 22218 10540 0 clknet_4_11_0_Clk
rlabel metal2 16974 14722 16974 14722 0 clknet_4_12_0_Clk
rlabel metal1 16606 20910 16606 20910 0 clknet_4_13_0_Clk
rlabel via1 19366 14909 19366 14909 0 clknet_4_14_0_Clk
rlabel metal1 20148 18258 20148 18258 0 clknet_4_15_0_Clk
rlabel metal1 2530 16116 2530 16116 0 clknet_4_1_0_Clk
rlabel metal1 6164 6766 6164 6766 0 clknet_4_2_0_Clk
rlabel metal1 7590 12886 7590 12886 0 clknet_4_3_0_Clk
rlabel metal1 7314 17646 7314 17646 0 clknet_4_4_0_Clk
rlabel metal1 4416 24174 4416 24174 0 clknet_4_5_0_Clk
rlabel metal1 13294 17204 13294 17204 0 clknet_4_6_0_Clk
rlabel metal2 9982 23936 9982 23936 0 clknet_4_7_0_Clk
rlabel metal2 14490 7038 14490 7038 0 clknet_4_8_0_Clk
rlabel metal1 13754 12750 13754 12750 0 clknet_4_9_0_Clk
rlabel metal1 8050 3468 8050 3468 0 fcounter\[0\]
rlabel metal1 11270 4046 11270 4046 0 fcounter\[1\]
rlabel metal2 9798 3536 9798 3536 0 fcounter\[2\]
rlabel metal2 5382 13396 5382 13396 0 memblk.FIFO\[0\]\[0\]
rlabel metal1 10948 18394 10948 18394 0 memblk.FIFO\[0\]\[10\]
rlabel metal1 11408 23834 11408 23834 0 memblk.FIFO\[0\]\[11\]
rlabel metal2 15318 18020 15318 18020 0 memblk.FIFO\[0\]\[12\]
rlabel metal1 15870 21658 15870 21658 0 memblk.FIFO\[0\]\[13\]
rlabel metal2 19274 24548 19274 24548 0 memblk.FIFO\[0\]\[14\]
rlabel metal2 15594 23868 15594 23868 0 memblk.FIFO\[0\]\[15\]
rlabel metal1 20194 21318 20194 21318 0 memblk.FIFO\[0\]\[16\]
rlabel metal1 19550 18292 19550 18292 0 memblk.FIFO\[0\]\[17\]
rlabel metal1 18446 11866 18446 11866 0 memblk.FIFO\[0\]\[18\]
rlabel metal2 21114 13702 21114 13702 0 memblk.FIFO\[0\]\[19\]
rlabel metal2 8786 10404 8786 10404 0 memblk.FIFO\[0\]\[1\]
rlabel metal2 23138 15028 23138 15028 0 memblk.FIFO\[0\]\[20\]
rlabel metal1 23552 17306 23552 17306 0 memblk.FIFO\[0\]\[21\]
rlabel metal1 18492 14586 18492 14586 0 memblk.FIFO\[0\]\[22\]
rlabel metal2 23598 10268 23598 10268 0 memblk.FIFO\[0\]\[23\]
rlabel metal1 19964 9146 19964 9146 0 memblk.FIFO\[0\]\[24\]
rlabel metal1 17434 6664 17434 6664 0 memblk.FIFO\[0\]\[25\]
rlabel metal1 22241 4046 22241 4046 0 memblk.FIFO\[0\]\[26\]
rlabel metal1 17388 4454 17388 4454 0 memblk.FIFO\[0\]\[27\]
rlabel metal1 22770 6324 22770 6324 0 memblk.FIFO\[0\]\[28\]
rlabel metal1 15824 10098 15824 10098 0 memblk.FIFO\[0\]\[29\]
rlabel metal1 5566 8466 5566 8466 0 memblk.FIFO\[0\]\[2\]
rlabel metal1 13846 14586 13846 14586 0 memblk.FIFO\[0\]\[30\]
rlabel metal1 11960 12954 11960 12954 0 memblk.FIFO\[0\]\[31\]
rlabel metal1 3082 10132 3082 10132 0 memblk.FIFO\[0\]\[3\]
rlabel metal1 8234 14858 8234 14858 0 memblk.FIFO\[0\]\[4\]
rlabel metal2 6302 16354 6302 16354 0 memblk.FIFO\[0\]\[5\]
rlabel metal1 11178 20978 11178 20978 0 memblk.FIFO\[0\]\[6\]
rlabel metal1 6486 23562 6486 23562 0 memblk.FIFO\[0\]\[7\]
rlabel metal2 7130 20604 7130 20604 0 memblk.FIFO\[0\]\[8\]
rlabel metal2 7130 19108 7130 19108 0 memblk.FIFO\[0\]\[9\]
rlabel metal2 4646 14076 4646 14076 0 memblk.FIFO\[1\]\[0\]
rlabel metal2 11362 17476 11362 17476 0 memblk.FIFO\[1\]\[10\]
rlabel metal1 11730 23698 11730 23698 0 memblk.FIFO\[1\]\[11\]
rlabel metal2 15410 17680 15410 17680 0 memblk.FIFO\[1\]\[12\]
rlabel metal1 15364 20570 15364 20570 0 memblk.FIFO\[1\]\[13\]
rlabel metal1 20332 23290 20332 23290 0 memblk.FIFO\[1\]\[14\]
rlabel metal1 15962 22950 15962 22950 0 memblk.FIFO\[1\]\[15\]
rlabel metal1 20516 21114 20516 21114 0 memblk.FIFO\[1\]\[16\]
rlabel metal1 19688 17306 19688 17306 0 memblk.FIFO\[1\]\[17\]
rlabel metal1 18400 12682 18400 12682 0 memblk.FIFO\[1\]\[18\]
rlabel metal1 23276 12410 23276 12410 0 memblk.FIFO\[1\]\[19\]
rlabel metal1 8418 10982 8418 10982 0 memblk.FIFO\[1\]\[1\]
rlabel metal1 23000 15470 23000 15470 0 memblk.FIFO\[1\]\[20\]
rlabel metal2 23138 18564 23138 18564 0 memblk.FIFO\[1\]\[21\]
rlabel metal1 18538 15538 18538 15538 0 memblk.FIFO\[1\]\[22\]
rlabel metal1 22402 10030 22402 10030 0 memblk.FIFO\[1\]\[23\]
rlabel metal1 19458 9452 19458 9452 0 memblk.FIFO\[1\]\[24\]
rlabel metal1 17572 5678 17572 5678 0 memblk.FIFO\[1\]\[25\]
rlabel metal1 19550 4114 19550 4114 0 memblk.FIFO\[1\]\[26\]
rlabel metal1 17756 3706 17756 3706 0 memblk.FIFO\[1\]\[27\]
rlabel metal1 20424 7514 20424 7514 0 memblk.FIFO\[1\]\[28\]
rlabel metal1 15686 11628 15686 11628 0 memblk.FIFO\[1\]\[29\]
rlabel metal2 5566 8126 5566 8126 0 memblk.FIFO\[1\]\[2\]
rlabel metal2 13938 14416 13938 14416 0 memblk.FIFO\[1\]\[30\]
rlabel metal2 12558 11628 12558 11628 0 memblk.FIFO\[1\]\[31\]
rlabel metal1 5152 10982 5152 10982 0 memblk.FIFO\[1\]\[3\]
rlabel metal1 7544 14586 7544 14586 0 memblk.FIFO\[1\]\[4\]
rlabel metal2 6486 16864 6486 16864 0 memblk.FIFO\[1\]\[5\]
rlabel metal1 12673 21454 12673 21454 0 memblk.FIFO\[1\]\[6\]
rlabel metal2 7038 23596 7038 23596 0 memblk.FIFO\[1\]\[7\]
rlabel metal2 7038 21216 7038 21216 0 memblk.FIFO\[1\]\[8\]
rlabel metal1 6992 18734 6992 18734 0 memblk.FIFO\[1\]\[9\]
rlabel metal1 3634 13396 3634 13396 0 memblk.FIFO\[2\]\[0\]
rlabel metal2 9706 16830 9706 16830 0 memblk.FIFO\[2\]\[10\]
rlabel metal1 10120 23494 10120 23494 0 memblk.FIFO\[2\]\[11\]
rlabel via1 14477 18258 14477 18258 0 memblk.FIFO\[2\]\[12\]
rlabel via1 15146 20978 15146 20978 0 memblk.FIFO\[2\]\[13\]
rlabel metal1 18308 23290 18308 23290 0 memblk.FIFO\[2\]\[14\]
rlabel metal1 14628 23290 14628 23290 0 memblk.FIFO\[2\]\[15\]
rlabel via1 18985 20434 18985 20434 0 memblk.FIFO\[2\]\[16\]
rlabel via1 18709 18190 18709 18190 0 memblk.FIFO\[2\]\[17\]
rlabel metal1 17651 12750 17651 12750 0 memblk.FIFO\[2\]\[18\]
rlabel metal1 21482 12614 21482 12614 0 memblk.FIFO\[2\]\[19\]
rlabel metal1 7314 10982 7314 10982 0 memblk.FIFO\[2\]\[1\]
rlabel metal1 21666 14484 21666 14484 0 memblk.FIFO\[2\]\[20\]
rlabel via1 22665 18258 22665 18258 0 memblk.FIFO\[2\]\[21\]
rlabel metal1 16836 16558 16836 16558 0 memblk.FIFO\[2\]\[22\]
rlabel metal1 21022 10778 21022 10778 0 memblk.FIFO\[2\]\[23\]
rlabel via1 18433 9486 18433 9486 0 memblk.FIFO\[2\]\[24\]
rlabel metal1 15686 5202 15686 5202 0 memblk.FIFO\[2\]\[25\]
rlabel via1 20390 4114 20390 4114 0 memblk.FIFO\[2\]\[26\]
rlabel metal1 16238 4012 16238 4012 0 memblk.FIFO\[2\]\[27\]
rlabel metal1 21436 6154 21436 6154 0 memblk.FIFO\[2\]\[28\]
rlabel metal1 14306 8806 14306 8806 0 memblk.FIFO\[2\]\[29\]
rlabel metal1 3818 7990 3818 7990 0 memblk.FIFO\[2\]\[2\]
rlabel metal1 11316 15130 11316 15130 0 memblk.FIFO\[2\]\[30\]
rlabel metal2 11454 11696 11454 11696 0 memblk.FIFO\[2\]\[31\]
rlabel metal2 3910 10064 3910 10064 0 memblk.FIFO\[2\]\[3\]
rlabel metal2 8418 13328 8418 13328 0 memblk.FIFO\[2\]\[4\]
rlabel metal1 4715 16626 4715 16626 0 memblk.FIFO\[2\]\[5\]
rlabel metal2 9338 20774 9338 20774 0 memblk.FIFO\[2\]\[6\]
rlabel metal1 5428 24310 5428 24310 0 memblk.FIFO\[2\]\[7\]
rlabel metal1 5819 20978 5819 20978 0 memblk.FIFO\[2\]\[8\]
rlabel metal2 5290 18700 5290 18700 0 memblk.FIFO\[2\]\[9\]
rlabel metal1 3542 14042 3542 14042 0 memblk.FIFO\[3\]\[0\]
rlabel metal1 9430 17714 9430 17714 0 memblk.FIFO\[3\]\[10\]
rlabel metal2 10074 22882 10074 22882 0 memblk.FIFO\[3\]\[11\]
rlabel metal1 14306 19278 14306 19278 0 memblk.FIFO\[3\]\[12\]
rlabel via1 15042 20893 15042 20893 0 memblk.FIFO\[3\]\[13\]
rlabel metal1 18998 23630 18998 23630 0 memblk.FIFO\[3\]\[14\]
rlabel metal1 14168 23834 14168 23834 0 memblk.FIFO\[3\]\[15\]
rlabel metal1 19182 21998 19182 21998 0 memblk.FIFO\[3\]\[16\]
rlabel metal1 17802 18632 17802 18632 0 memblk.FIFO\[3\]\[17\]
rlabel metal1 16376 13294 16376 13294 0 memblk.FIFO\[3\]\[18\]
rlabel metal1 21344 13838 21344 13838 0 memblk.FIFO\[3\]\[19\]
rlabel metal2 5658 10404 5658 10404 0 memblk.FIFO\[3\]\[1\]
rlabel metal1 21114 16014 21114 16014 0 memblk.FIFO\[3\]\[20\]
rlabel metal1 22724 19278 22724 19278 0 memblk.FIFO\[3\]\[21\]
rlabel metal2 17066 14994 17066 14994 0 memblk.FIFO\[3\]\[22\]
rlabel metal1 23414 11254 23414 11254 0 memblk.FIFO\[3\]\[23\]
rlabel metal1 18446 10132 18446 10132 0 memblk.FIFO\[3\]\[24\]
rlabel metal2 15502 6732 15502 6732 0 memblk.FIFO\[3\]\[25\]
rlabel metal1 19964 4590 19964 4590 0 memblk.FIFO\[3\]\[26\]
rlabel metal1 15134 4046 15134 4046 0 memblk.FIFO\[3\]\[27\]
rlabel metal2 20102 6868 20102 6868 0 memblk.FIFO\[3\]\[28\]
rlabel via1 15042 10115 15042 10115 0 memblk.FIFO\[3\]\[29\]
rlabel metal1 3818 8942 3818 8942 0 memblk.FIFO\[3\]\[2\]
rlabel metal2 13018 15504 13018 15504 0 memblk.FIFO\[3\]\[30\]
rlabel metal1 11178 12750 11178 12750 0 memblk.FIFO\[3\]\[31\]
rlabel metal1 3450 11662 3450 11662 0 memblk.FIFO\[3\]\[3\]
rlabel metal1 7222 13498 7222 13498 0 memblk.FIFO\[3\]\[4\]
rlabel metal1 5658 16626 5658 16626 0 memblk.FIFO\[3\]\[5\]
rlabel metal2 10350 21658 10350 21658 0 memblk.FIFO\[3\]\[6\]
rlabel metal2 6118 23324 6118 23324 0 memblk.FIFO\[3\]\[7\]
rlabel metal1 5382 21318 5382 21318 0 memblk.FIFO\[3\]\[8\]
rlabel metal1 6026 19312 6026 19312 0 memblk.FIFO\[3\]\[9\]
rlabel metal1 13386 13226 13386 13226 0 memblk.rd_addr\[0\]
rlabel metal1 16284 10710 16284 10710 0 memblk.rd_addr\[1\]
rlabel metal2 13294 5848 13294 5848 0 memblk.wr_addr\[0\]
rlabel metal1 12926 7888 12926 7888 0 memblk.wr_addr\[1\]
rlabel metal2 2714 14620 2714 14620 0 net1
rlabel metal2 18722 11934 18722 11934 0 net10
rlabel metal1 21712 11050 21712 11050 0 net100
rlabel metal1 5244 18394 5244 18394 0 net101
rlabel metal1 17710 22746 17710 22746 0 net102
rlabel metal1 4692 18666 4692 18666 0 net103
rlabel metal2 11546 17408 11546 17408 0 net104
rlabel metal2 23046 10608 23046 10608 0 net105
rlabel metal1 10534 18666 10534 18666 0 net106
rlabel metal2 9430 23868 9430 23868 0 net107
rlabel metal2 17158 9248 17158 9248 0 net108
rlabel metal2 15778 10064 15778 10064 0 net109
rlabel metal1 22218 11662 22218 11662 0 net11
rlabel metal1 8004 15130 8004 15130 0 net110
rlabel metal2 16054 18496 16054 18496 0 net111
rlabel metal2 2622 13090 2622 13090 0 net112
rlabel metal1 21528 10778 21528 10778 0 net113
rlabel metal1 8970 17170 8970 17170 0 net114
rlabel metal1 6946 20366 6946 20366 0 net115
rlabel metal2 18538 21386 18538 21386 0 net116
rlabel metal1 17940 7922 17940 7922 0 net117
rlabel metal1 9384 22746 9384 22746 0 net118
rlabel metal1 16192 14314 16192 14314 0 net119
rlabel metal2 9338 10166 9338 10166 0 net12
rlabel metal2 16974 3842 16974 3842 0 net120
rlabel metal2 5750 24242 5750 24242 0 net121
rlabel metal1 3082 9554 3082 9554 0 net122
rlabel metal2 21022 14756 21022 14756 0 net123
rlabel metal2 7866 13056 7866 13056 0 net124
rlabel metal2 14490 21760 14490 21760 0 net125
rlabel metal1 20562 23698 20562 23698 0 net126
rlabel metal1 18998 4522 18998 4522 0 net127
rlabel metal1 5796 9146 5796 9146 0 net128
rlabel metal2 6394 8704 6394 8704 0 net129
rlabel metal1 20976 14994 20976 14994 0 net13
rlabel metal2 18354 23834 18354 23834 0 net130
rlabel metal1 4094 15130 4094 15130 0 net131
rlabel metal1 7176 18326 7176 18326 0 net132
rlabel metal1 8142 9554 8142 9554 0 net133
rlabel metal2 4462 16320 4462 16320 0 net134
rlabel metal2 18906 8976 18906 8976 0 net135
rlabel metal2 19274 11968 19274 11968 0 net136
rlabel metal2 19734 8092 19734 8092 0 net137
rlabel metal2 15870 23494 15870 23494 0 net138
rlabel metal2 9430 19584 9430 19584 0 net139
rlabel metal1 21574 17544 21574 17544 0 net14
rlabel metal1 17894 16082 17894 16082 0 net140
rlabel metal1 22678 16490 22678 16490 0 net141
rlabel metal2 10994 15708 10994 15708 0 net142
rlabel metal2 14582 16830 14582 16830 0 net143
rlabel metal1 9430 14450 9430 14450 0 net144
rlabel metal1 13616 19346 13616 19346 0 net145
rlabel metal2 15318 5984 15318 5984 0 net146
rlabel metal2 13846 9248 13846 9248 0 net147
rlabel metal1 6486 7718 6486 7718 0 net148
rlabel metal1 12190 21522 12190 21522 0 net149
rlabel metal2 18814 15232 18814 15232 0 net15
rlabel metal1 19090 14586 19090 14586 0 net150
rlabel metal1 22540 11730 22540 11730 0 net151
rlabel metal1 18814 16626 18814 16626 0 net152
rlabel metal2 6854 22848 6854 22848 0 net153
rlabel metal1 20930 7786 20930 7786 0 net154
rlabel metal2 15410 3536 15410 3536 0 net155
rlabel metal1 10626 19924 10626 19924 0 net156
rlabel metal2 15962 16320 15962 16320 0 net157
rlabel metal2 19734 18972 19734 18972 0 net158
rlabel metal1 20286 5134 20286 5134 0 net159
rlabel metal2 22034 9316 22034 9316 0 net16
rlabel metal2 21390 13532 21390 13532 0 net160
rlabel metal1 15042 19686 15042 19686 0 net161
rlabel metal1 7038 21522 7038 21522 0 net162
rlabel metal1 14674 14586 14674 14586 0 net163
rlabel metal1 21850 17680 21850 17680 0 net164
rlabel metal1 6118 17170 6118 17170 0 net165
rlabel metal1 21114 3094 21114 3094 0 net166
rlabel metal1 14352 22678 14352 22678 0 net167
rlabel metal1 23874 15674 23874 15674 0 net168
rlabel metal1 11776 13158 11776 13158 0 net169
rlabel metal1 19780 7854 19780 7854 0 net17
rlabel metal1 11132 24786 11132 24786 0 net170
rlabel metal1 17894 19686 17894 19686 0 net171
rlabel metal1 22402 13838 22402 13838 0 net172
rlabel metal1 11270 22746 11270 22746 0 net173
rlabel metal2 16514 11968 16514 11968 0 net174
rlabel metal1 15318 22610 15318 22610 0 net175
rlabel metal1 5382 13906 5382 13906 0 net176
rlabel metal2 9430 11152 9430 11152 0 net177
rlabel metal1 7038 16082 7038 16082 0 net178
rlabel metal2 19734 3264 19734 3264 0 net179
rlabel metal1 16606 2618 16606 2618 0 net18
rlabel metal2 21206 21148 21206 21148 0 net180
rlabel metal1 17342 4250 17342 4250 0 net181
rlabel metal1 14950 11730 14950 11730 0 net182
rlabel metal1 5382 21862 5382 21862 0 net183
rlabel metal2 21114 16932 21114 16932 0 net184
rlabel metal2 18262 18156 18262 18156 0 net185
rlabel metal1 3358 6970 3358 6970 0 net186
rlabel metal1 4876 22610 4876 22610 0 net187
rlabel metal1 10626 11050 10626 11050 0 net188
rlabel metal1 17342 7378 17342 7378 0 net189
rlabel metal1 19688 2618 19688 2618 0 net19
rlabel metal2 20700 12852 20700 12852 0 net190
rlabel metal2 6854 10574 6854 10574 0 net191
rlabel metal1 17250 9690 17250 9690 0 net192
rlabel metal1 18906 24242 18906 24242 0 net193
rlabel metal2 15686 21216 15686 21216 0 net194
rlabel metal1 4370 11730 4370 11730 0 net195
rlabel metal2 18630 21760 18630 21760 0 net196
rlabel metal1 13754 13294 13754 13294 0 net197
rlabel metal1 20516 7446 20516 7446 0 net198
rlabel metal1 4370 9622 4370 9622 0 net199
rlabel metal1 8464 24582 8464 24582 0 net2
rlabel metal1 15548 2618 15548 2618 0 net20
rlabel metal1 17342 5338 17342 5338 0 net200
rlabel metal1 17940 11050 17940 11050 0 net201
rlabel metal1 11454 11322 11454 11322 0 net202
rlabel metal2 22218 5950 22218 5950 0 net203
rlabel metal1 12236 7378 12236 7378 0 net204
rlabel metal1 23506 6188 23506 6188 0 net21
rlabel metal1 14444 2618 14444 2618 0 net22
rlabel metal2 5014 8296 5014 8296 0 net23
rlabel metal1 14076 15062 14076 15062 0 net24
rlabel metal1 10258 12750 10258 12750 0 net25
rlabel metal1 2185 11866 2185 11866 0 net26
rlabel metal1 1610 15368 1610 15368 0 net27
rlabel metal1 4370 15980 4370 15980 0 net28
rlabel metal1 9108 21998 9108 21998 0 net29
rlabel metal1 9430 22950 9430 22950 0 net3
rlabel metal1 6302 23698 6302 23698 0 net30
rlabel metal1 4968 24650 4968 24650 0 net31
rlabel metal1 2185 18870 2185 18870 0 net32
rlabel metal1 10764 3978 10764 3978 0 net33
rlabel metal1 12236 2550 12236 2550 0 net34
rlabel metal2 8050 3094 8050 3094 0 net35
rlabel metal1 6670 2618 6670 2618 0 net36
rlabel metal1 1840 12818 1840 12818 0 net37
rlabel metal2 11592 23596 11592 23596 0 net38
rlabel metal2 12466 24582 12466 24582 0 net39
rlabel metal1 13386 19482 13386 19482 0 net4
rlabel metal1 15272 19482 15272 19482 0 net40
rlabel metal1 16146 21114 16146 21114 0 net41
rlabel metal1 20976 23834 20976 23834 0 net42
rlabel metal2 16238 24582 16238 24582 0 net43
rlabel metal1 20930 20570 20930 20570 0 net44
rlabel metal2 20010 18530 20010 18530 0 net45
rlabel metal1 23322 12206 23322 12206 0 net46
rlabel metal1 22770 10778 22770 10778 0 net47
rlabel metal1 2070 11220 2070 11220 0 net48
rlabel metal1 22218 17306 22218 17306 0 net49
rlabel metal2 14766 20128 14766 20128 0 net5
rlabel metal1 23276 19346 23276 19346 0 net50
rlabel metal1 19550 15674 19550 15674 0 net51
rlabel metal1 22908 9146 22908 9146 0 net52
rlabel metal1 22678 9656 22678 9656 0 net53
rlabel metal1 18170 2346 18170 2346 0 net54
rlabel metal2 21942 2890 21942 2890 0 net55
rlabel metal1 17388 2414 17388 2414 0 net56
rlabel metal1 23138 7378 23138 7378 0 net57
rlabel metal1 14812 2414 14812 2414 0 net58
rlabel metal1 3450 8432 3450 8432 0 net59
rlabel metal1 19182 24106 19182 24106 0 net6
rlabel metal2 15870 14144 15870 14144 0 net60
rlabel metal1 12788 2414 12788 2414 0 net61
rlabel metal2 1702 11356 1702 11356 0 net62
rlabel metal1 1702 14484 1702 14484 0 net63
rlabel metal1 1702 16490 1702 16490 0 net64
rlabel metal1 11776 24106 11776 24106 0 net65
rlabel metal2 7866 23970 7866 23970 0 net66
rlabel metal1 7268 24786 7268 24786 0 net67
rlabel metal1 1702 19414 1702 19414 0 net68
rlabel metal1 7590 2448 7590 2448 0 net69
rlabel metal2 14674 22882 14674 22882 0 net7
rlabel metal1 6716 2414 6716 2414 0 net70
rlabel metal1 8648 2414 8648 2414 0 net71
rlabel metal1 9936 2482 9936 2482 0 net72
rlabel metal1 7981 6630 7981 6630 0 net73
rlabel metal2 11546 8364 11546 8364 0 net74
rlabel metal1 7682 3638 7682 3638 0 net75
rlabel metal1 13846 24174 13846 24174 0 net76
rlabel metal1 14766 3502 14766 3502 0 net77
rlabel metal1 4922 22746 4922 22746 0 net78
rlabel metal1 10488 12818 10488 12818 0 net79
rlabel metal2 18630 20298 18630 20298 0 net8
rlabel metal2 2806 11322 2806 11322 0 net80
rlabel metal1 16008 13226 16008 13226 0 net81
rlabel metal1 3450 8874 3450 8874 0 net82
rlabel metal2 6946 14144 6946 14144 0 net83
rlabel metal1 20700 16082 20700 16082 0 net84
rlabel metal1 4416 20910 4416 20910 0 net85
rlabel metal1 2852 14382 2852 14382 0 net86
rlabel metal1 6992 18394 6992 18394 0 net87
rlabel metal2 13570 21760 13570 21760 0 net88
rlabel metal1 15870 6426 15870 6426 0 net89
rlabel metal1 19780 18734 19780 18734 0 net9
rlabel metal1 4462 14246 4462 14246 0 net90
rlabel metal1 22494 9554 22494 9554 0 net91
rlabel metal1 20884 12954 20884 12954 0 net92
rlabel metal2 22126 18972 22126 18972 0 net93
rlabel metal2 11730 15674 11730 15674 0 net94
rlabel metal1 13800 18598 13800 18598 0 net95
rlabel metal2 8786 18496 8786 18496 0 net96
rlabel metal1 9568 21930 9568 21930 0 net97
rlabel metal1 17710 17306 17710 17306 0 net98
rlabel metal1 19228 6766 19228 6766 0 net99
<< properties >>
string FIXED_BBOX 0 0 25180 27324
<< end >>
