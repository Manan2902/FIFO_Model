VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FIFO_Model
  CLASS BLOCK ;
  FOREIGN FIFO_Model ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.900 BY 136.620 ;
  PIN Clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END Clk
  PIN Data_In[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.000 68.640 ;
    END
  END Data_In[0]
  PIN Data_In[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 134.620 42.230 136.620 ;
    END
  END Data_In[10]
  PIN Data_In[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 134.620 48.670 136.620 ;
    END
  END Data_In[11]
  PIN Data_In[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 134.620 64.770 136.620 ;
    END
  END Data_In[12]
  PIN Data_In[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 134.620 71.210 136.620 ;
    END
  END Data_In[13]
  PIN Data_In[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 134.620 93.750 136.620 ;
    END
  END Data_In[14]
  PIN Data_In[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 134.620 67.990 136.620 ;
    END
  END Data_In[15]
  PIN Data_In[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 134.620 96.970 136.620 ;
    END
  END Data_In[16]
  PIN Data_In[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 98.640 125.900 99.240 ;
    END
  END Data_In[17]
  PIN Data_In[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 57.840 125.900 58.440 ;
    END
  END Data_In[18]
  PIN Data_In[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 68.040 125.900 68.640 ;
    END
  END Data_In[19]
  PIN Data_In[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.000 48.240 ;
    END
  END Data_In[1]
  PIN Data_In[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 74.840 125.900 75.440 ;
    END
  END Data_In[20]
  PIN Data_In[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 88.440 125.900 89.040 ;
    END
  END Data_In[21]
  PIN Data_In[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 85.040 125.900 85.640 ;
    END
  END Data_In[22]
  PIN Data_In[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 54.440 125.900 55.040 ;
    END
  END Data_In[23]
  PIN Data_In[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 44.240 125.900 44.840 ;
    END
  END Data_In[24]
  PIN Data_In[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.000 ;
    END
  END Data_In[25]
  PIN Data_In[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.000 ;
    END
  END Data_In[26]
  PIN Data_In[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.000 ;
    END
  END Data_In[27]
  PIN Data_In[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 30.640 125.900 31.240 ;
    END
  END Data_In[28]
  PIN Data_In[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 2.000 ;
    END
  END Data_In[29]
  PIN Data_In[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.000 44.840 ;
    END
  END Data_In[2]
  PIN Data_In[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 134.620 61.550 136.620 ;
    END
  END Data_In[30]
  PIN Data_In[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.000 61.840 ;
    END
  END Data_In[31]
  PIN Data_In[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.000 58.440 ;
    END
  END Data_In[3]
  PIN Data_In[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.000 75.440 ;
    END
  END Data_In[4]
  PIN Data_In[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END Data_In[5]
  PIN Data_In[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 134.620 45.450 136.620 ;
    END
  END Data_In[6]
  PIN Data_In[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 134.620 29.350 136.620 ;
    END
  END Data_In[7]
  PIN Data_In[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 134.620 26.130 136.620 ;
    END
  END Data_In[8]
  PIN Data_In[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.000 92.440 ;
    END
  END Data_In[9]
  PIN FClrN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.000 ;
    END
  END FClrN
  PIN FInN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.000 ;
    END
  END FInN
  PIN FOutN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.000 ;
    END
  END FOutN
  PIN F_Data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.000 65.240 ;
    END
  END F_Data[0]
  PIN F_Data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 134.620 51.890 136.620 ;
    END
  END F_Data[10]
  PIN F_Data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.050 134.620 58.330 136.620 ;
    END
  END F_Data[11]
  PIN F_Data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 134.620 74.430 136.620 ;
    END
  END F_Data[12]
  PIN F_Data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 134.620 80.870 136.620 ;
    END
  END F_Data[13]
  PIN F_Data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.910 134.620 100.190 136.620 ;
    END
  END F_Data[14]
  PIN F_Data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 134.620 77.650 136.620 ;
    END
  END F_Data[15]
  PIN F_Data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 105.440 125.900 106.040 ;
    END
  END F_Data[16]
  PIN F_Data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 91.840 125.900 92.440 ;
    END
  END F_Data[17]
  PIN F_Data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 61.240 125.900 61.840 ;
    END
  END F_Data[18]
  PIN F_Data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 64.640 125.900 65.240 ;
    END
  END F_Data[19]
  PIN F_Data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 2.000 51.640 ;
    END
  END F_Data[1]
  PIN F_Data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 81.640 125.900 82.240 ;
    END
  END F_Data[20]
  PIN F_Data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 95.240 125.900 95.840 ;
    END
  END F_Data[21]
  PIN F_Data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 78.240 125.900 78.840 ;
    END
  END F_Data[22]
  PIN F_Data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 51.040 125.900 51.640 ;
    END
  END F_Data[23]
  PIN F_Data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 47.640 125.900 48.240 ;
    END
  END F_Data[24]
  PIN F_Data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.000 ;
    END
  END F_Data[25]
  PIN F_Data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 2.000 ;
    END
  END F_Data[26]
  PIN F_Data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.000 ;
    END
  END F_Data[27]
  PIN F_Data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 34.040 125.900 34.640 ;
    END
  END F_Data[28]
  PIN F_Data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 2.000 ;
    END
  END F_Data[29]
  PIN F_Data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END F_Data[2]
  PIN F_Data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 123.900 71.440 125.900 72.040 ;
    END
  END F_Data[30]
  PIN F_Data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.000 ;
    END
  END F_Data[31]
  PIN F_Data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 2.000 55.040 ;
    END
  END F_Data[3]
  PIN F_Data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.000 72.040 ;
    END
  END F_Data[4]
  PIN F_Data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.000 82.240 ;
    END
  END F_Data[5]
  PIN F_Data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 134.620 55.110 136.620 ;
    END
  END F_Data[6]
  PIN F_Data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 134.620 32.570 136.620 ;
    END
  END F_Data[7]
  PIN F_Data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 134.620 35.790 136.620 ;
    END
  END F_Data[8]
  PIN F_Data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.000 95.840 ;
    END
  END F_Data[9]
  PIN F_EmptyN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.000 ;
    END
  END F_EmptyN
  PIN F_FirstN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.000 ;
    END
  END F_FirstN
  PIN F_FullN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.000 ;
    END
  END F_FullN
  PIN F_LastN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 2.000 ;
    END
  END F_LastN
  PIN F_SLastN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.000 ;
    END
  END F_SLastN
  PIN RstN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.000 ;
    END
  END RstN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.220 10.640 15.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.220 10.640 30.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.220 10.640 45.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.220 10.640 60.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.220 10.640 75.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.220 10.640 90.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.220 10.640 105.820 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.220 10.640 120.820 125.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.720 10.640 8.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.720 10.640 23.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.720 10.640 38.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.720 10.640 53.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.720 10.640 68.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.720 10.640 83.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.720 10.640 98.320 125.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.720 10.640 113.320 125.360 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 120.250 125.205 ;
      LAYER li1 ;
        RECT 5.520 10.795 120.060 125.205 ;
      LAYER met1 ;
        RECT 1.910 10.640 121.830 125.360 ;
      LAYER met2 ;
        RECT 1.930 134.340 25.570 135.050 ;
        RECT 26.410 134.340 28.790 135.050 ;
        RECT 29.630 134.340 32.010 135.050 ;
        RECT 32.850 134.340 35.230 135.050 ;
        RECT 36.070 134.340 41.670 135.050 ;
        RECT 42.510 134.340 44.890 135.050 ;
        RECT 45.730 134.340 48.110 135.050 ;
        RECT 48.950 134.340 51.330 135.050 ;
        RECT 52.170 134.340 54.550 135.050 ;
        RECT 55.390 134.340 57.770 135.050 ;
        RECT 58.610 134.340 60.990 135.050 ;
        RECT 61.830 134.340 64.210 135.050 ;
        RECT 65.050 134.340 67.430 135.050 ;
        RECT 68.270 134.340 70.650 135.050 ;
        RECT 71.490 134.340 73.870 135.050 ;
        RECT 74.710 134.340 77.090 135.050 ;
        RECT 77.930 134.340 80.310 135.050 ;
        RECT 81.150 134.340 93.190 135.050 ;
        RECT 94.030 134.340 96.410 135.050 ;
        RECT 97.250 134.340 99.630 135.050 ;
        RECT 100.470 134.340 121.810 135.050 ;
        RECT 1.930 2.280 121.810 134.340 ;
        RECT 1.930 2.000 28.790 2.280 ;
        RECT 29.630 2.000 32.010 2.280 ;
        RECT 32.850 2.000 35.230 2.280 ;
        RECT 36.070 2.000 38.450 2.280 ;
        RECT 39.290 2.000 41.670 2.280 ;
        RECT 42.510 2.000 44.890 2.280 ;
        RECT 45.730 2.000 48.110 2.280 ;
        RECT 48.950 2.000 51.330 2.280 ;
        RECT 52.170 2.000 57.770 2.280 ;
        RECT 58.610 2.000 60.990 2.280 ;
        RECT 61.830 2.000 70.650 2.280 ;
        RECT 71.490 2.000 73.870 2.280 ;
        RECT 74.710 2.000 77.090 2.280 ;
        RECT 77.930 2.000 80.310 2.280 ;
        RECT 81.150 2.000 83.530 2.280 ;
        RECT 84.370 2.000 86.750 2.280 ;
        RECT 87.590 2.000 96.410 2.280 ;
        RECT 97.250 2.000 106.070 2.280 ;
        RECT 106.910 2.000 121.810 2.280 ;
      LAYER met3 ;
        RECT 2.000 116.640 123.900 125.285 ;
        RECT 2.400 115.240 123.900 116.640 ;
        RECT 2.000 106.440 123.900 115.240 ;
        RECT 2.000 105.040 123.500 106.440 ;
        RECT 2.000 99.640 123.900 105.040 ;
        RECT 2.000 98.240 123.500 99.640 ;
        RECT 2.000 96.240 123.900 98.240 ;
        RECT 2.400 94.840 123.500 96.240 ;
        RECT 2.000 92.840 123.900 94.840 ;
        RECT 2.400 91.440 123.500 92.840 ;
        RECT 2.000 89.440 123.900 91.440 ;
        RECT 2.000 88.040 123.500 89.440 ;
        RECT 2.000 86.040 123.900 88.040 ;
        RECT 2.000 84.640 123.500 86.040 ;
        RECT 2.000 82.640 123.900 84.640 ;
        RECT 2.400 81.240 123.500 82.640 ;
        RECT 2.000 79.240 123.900 81.240 ;
        RECT 2.400 77.840 123.500 79.240 ;
        RECT 2.000 75.840 123.900 77.840 ;
        RECT 2.400 74.440 123.500 75.840 ;
        RECT 2.000 72.440 123.900 74.440 ;
        RECT 2.400 71.040 123.500 72.440 ;
        RECT 2.000 69.040 123.900 71.040 ;
        RECT 2.400 67.640 123.500 69.040 ;
        RECT 2.000 65.640 123.900 67.640 ;
        RECT 2.400 64.240 123.500 65.640 ;
        RECT 2.000 62.240 123.900 64.240 ;
        RECT 2.400 60.840 123.500 62.240 ;
        RECT 2.000 58.840 123.900 60.840 ;
        RECT 2.400 57.440 123.500 58.840 ;
        RECT 2.000 55.440 123.900 57.440 ;
        RECT 2.400 54.040 123.500 55.440 ;
        RECT 2.000 52.040 123.900 54.040 ;
        RECT 2.400 50.640 123.500 52.040 ;
        RECT 2.000 48.640 123.900 50.640 ;
        RECT 2.400 47.240 123.500 48.640 ;
        RECT 2.000 45.240 123.900 47.240 ;
        RECT 2.400 43.840 123.500 45.240 ;
        RECT 2.000 41.840 123.900 43.840 ;
        RECT 2.400 40.440 123.900 41.840 ;
        RECT 2.000 35.040 123.900 40.440 ;
        RECT 2.000 33.640 123.500 35.040 ;
        RECT 2.000 31.640 123.900 33.640 ;
        RECT 2.000 30.240 123.500 31.640 ;
        RECT 2.000 10.715 123.900 30.240 ;
      LAYER met4 ;
        RECT 16.855 55.255 21.320 116.105 ;
        RECT 23.720 55.255 28.820 116.105 ;
        RECT 31.220 55.255 36.320 116.105 ;
        RECT 38.720 55.255 43.820 116.105 ;
        RECT 46.220 55.255 51.320 116.105 ;
        RECT 53.720 55.255 58.820 116.105 ;
        RECT 61.220 55.255 66.320 116.105 ;
        RECT 68.720 55.255 73.820 116.105 ;
        RECT 76.220 55.255 81.320 116.105 ;
        RECT 83.720 55.255 88.820 116.105 ;
        RECT 91.220 55.255 96.320 116.105 ;
        RECT 98.720 55.255 103.820 116.105 ;
        RECT 106.220 55.255 111.025 116.105 ;
  END
END FIFO_Model
END LIBRARY

