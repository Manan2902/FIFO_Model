module FIFO_Model (Clk,
    FClrN,
    FInN,
    FOutN,
    F_EmptyN,
    F_FirstN,
    F_FullN,
    F_LastN,
    F_SLastN,
    RstN,
    Data_In,
    F_Data);
 input Clk;
 input FClrN;
 input FInN;
 input FOutN;
 output F_EmptyN;
 output F_FirstN;
 output F_FullN;
 output F_LastN;
 output F_SLastN;
 input RstN;
 input [31:0] Data_In;
 output [31:0] F_Data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire \fcounter[0] ;
 wire \fcounter[1] ;
 wire \fcounter[2] ;
 wire \memblk.FIFO[0][0] ;
 wire \memblk.FIFO[0][10] ;
 wire \memblk.FIFO[0][11] ;
 wire \memblk.FIFO[0][12] ;
 wire \memblk.FIFO[0][13] ;
 wire \memblk.FIFO[0][14] ;
 wire \memblk.FIFO[0][15] ;
 wire \memblk.FIFO[0][16] ;
 wire \memblk.FIFO[0][17] ;
 wire \memblk.FIFO[0][18] ;
 wire \memblk.FIFO[0][19] ;
 wire \memblk.FIFO[0][1] ;
 wire \memblk.FIFO[0][20] ;
 wire \memblk.FIFO[0][21] ;
 wire \memblk.FIFO[0][22] ;
 wire \memblk.FIFO[0][23] ;
 wire \memblk.FIFO[0][24] ;
 wire \memblk.FIFO[0][25] ;
 wire \memblk.FIFO[0][26] ;
 wire \memblk.FIFO[0][27] ;
 wire \memblk.FIFO[0][28] ;
 wire \memblk.FIFO[0][29] ;
 wire \memblk.FIFO[0][2] ;
 wire \memblk.FIFO[0][30] ;
 wire \memblk.FIFO[0][31] ;
 wire \memblk.FIFO[0][3] ;
 wire \memblk.FIFO[0][4] ;
 wire \memblk.FIFO[0][5] ;
 wire \memblk.FIFO[0][6] ;
 wire \memblk.FIFO[0][7] ;
 wire \memblk.FIFO[0][8] ;
 wire \memblk.FIFO[0][9] ;
 wire \memblk.FIFO[1][0] ;
 wire \memblk.FIFO[1][10] ;
 wire \memblk.FIFO[1][11] ;
 wire \memblk.FIFO[1][12] ;
 wire \memblk.FIFO[1][13] ;
 wire \memblk.FIFO[1][14] ;
 wire \memblk.FIFO[1][15] ;
 wire \memblk.FIFO[1][16] ;
 wire \memblk.FIFO[1][17] ;
 wire \memblk.FIFO[1][18] ;
 wire \memblk.FIFO[1][19] ;
 wire \memblk.FIFO[1][1] ;
 wire \memblk.FIFO[1][20] ;
 wire \memblk.FIFO[1][21] ;
 wire \memblk.FIFO[1][22] ;
 wire \memblk.FIFO[1][23] ;
 wire \memblk.FIFO[1][24] ;
 wire \memblk.FIFO[1][25] ;
 wire \memblk.FIFO[1][26] ;
 wire \memblk.FIFO[1][27] ;
 wire \memblk.FIFO[1][28] ;
 wire \memblk.FIFO[1][29] ;
 wire \memblk.FIFO[1][2] ;
 wire \memblk.FIFO[1][30] ;
 wire \memblk.FIFO[1][31] ;
 wire \memblk.FIFO[1][3] ;
 wire \memblk.FIFO[1][4] ;
 wire \memblk.FIFO[1][5] ;
 wire \memblk.FIFO[1][6] ;
 wire \memblk.FIFO[1][7] ;
 wire \memblk.FIFO[1][8] ;
 wire \memblk.FIFO[1][9] ;
 wire \memblk.FIFO[2][0] ;
 wire \memblk.FIFO[2][10] ;
 wire \memblk.FIFO[2][11] ;
 wire \memblk.FIFO[2][12] ;
 wire \memblk.FIFO[2][13] ;
 wire \memblk.FIFO[2][14] ;
 wire \memblk.FIFO[2][15] ;
 wire \memblk.FIFO[2][16] ;
 wire \memblk.FIFO[2][17] ;
 wire \memblk.FIFO[2][18] ;
 wire \memblk.FIFO[2][19] ;
 wire \memblk.FIFO[2][1] ;
 wire \memblk.FIFO[2][20] ;
 wire \memblk.FIFO[2][21] ;
 wire \memblk.FIFO[2][22] ;
 wire \memblk.FIFO[2][23] ;
 wire \memblk.FIFO[2][24] ;
 wire \memblk.FIFO[2][25] ;
 wire \memblk.FIFO[2][26] ;
 wire \memblk.FIFO[2][27] ;
 wire \memblk.FIFO[2][28] ;
 wire \memblk.FIFO[2][29] ;
 wire \memblk.FIFO[2][2] ;
 wire \memblk.FIFO[2][30] ;
 wire \memblk.FIFO[2][31] ;
 wire \memblk.FIFO[2][3] ;
 wire \memblk.FIFO[2][4] ;
 wire \memblk.FIFO[2][5] ;
 wire \memblk.FIFO[2][6] ;
 wire \memblk.FIFO[2][7] ;
 wire \memblk.FIFO[2][8] ;
 wire \memblk.FIFO[2][9] ;
 wire \memblk.FIFO[3][0] ;
 wire \memblk.FIFO[3][10] ;
 wire \memblk.FIFO[3][11] ;
 wire \memblk.FIFO[3][12] ;
 wire \memblk.FIFO[3][13] ;
 wire \memblk.FIFO[3][14] ;
 wire \memblk.FIFO[3][15] ;
 wire \memblk.FIFO[3][16] ;
 wire \memblk.FIFO[3][17] ;
 wire \memblk.FIFO[3][18] ;
 wire \memblk.FIFO[3][19] ;
 wire \memblk.FIFO[3][1] ;
 wire \memblk.FIFO[3][20] ;
 wire \memblk.FIFO[3][21] ;
 wire \memblk.FIFO[3][22] ;
 wire \memblk.FIFO[3][23] ;
 wire \memblk.FIFO[3][24] ;
 wire \memblk.FIFO[3][25] ;
 wire \memblk.FIFO[3][26] ;
 wire \memblk.FIFO[3][27] ;
 wire \memblk.FIFO[3][28] ;
 wire \memblk.FIFO[3][29] ;
 wire \memblk.FIFO[3][2] ;
 wire \memblk.FIFO[3][30] ;
 wire \memblk.FIFO[3][31] ;
 wire \memblk.FIFO[3][3] ;
 wire \memblk.FIFO[3][4] ;
 wire \memblk.FIFO[3][5] ;
 wire \memblk.FIFO[3][6] ;
 wire \memblk.FIFO[3][7] ;
 wire \memblk.FIFO[3][8] ;
 wire \memblk.FIFO[3][9] ;
 wire \memblk.rd_addr[0] ;
 wire \memblk.rd_addr[1] ;
 wire \memblk.wr_addr[0] ;
 wire \memblk.wr_addr[1] ;

 sky130_fd_sc_hd__buf_2 _389_ (.A(\memblk.rd_addr[0] ),
    .X(_140_));
 sky130_fd_sc_hd__buf_2 _390_ (.A(_140_),
    .X(_141_));
 sky130_fd_sc_hd__buf_1 _391_ (.A(\memblk.rd_addr[1] ),
    .X(_142_));
 sky130_fd_sc_hd__buf_1 _392_ (.A(_142_),
    .X(_143_));
 sky130_fd_sc_hd__mux4_2 _393_ (.A0(\memblk.FIFO[0][0] ),
    .A1(\memblk.FIFO[1][0] ),
    .A2(\memblk.FIFO[2][0] ),
    .A3(\memblk.FIFO[3][0] ),
    .S0(_141_),
    .S1(_143_),
    .X(_144_));
 sky130_fd_sc_hd__buf_1 _394_ (.A(_144_),
    .X(F_Data[0]));
 sky130_fd_sc_hd__mux4_2 _395_ (.A0(\memblk.FIFO[0][1] ),
    .A1(\memblk.FIFO[1][1] ),
    .A2(\memblk.FIFO[2][1] ),
    .A3(\memblk.FIFO[3][1] ),
    .S0(_141_),
    .S1(_143_),
    .X(_145_));
 sky130_fd_sc_hd__buf_1 _396_ (.A(_145_),
    .X(F_Data[1]));
 sky130_fd_sc_hd__mux4_2 _397_ (.A0(\memblk.FIFO[0][2] ),
    .A1(\memblk.FIFO[1][2] ),
    .A2(\memblk.FIFO[2][2] ),
    .A3(\memblk.FIFO[3][2] ),
    .S0(_141_),
    .S1(_143_),
    .X(_146_));
 sky130_fd_sc_hd__buf_1 _398_ (.A(_146_),
    .X(F_Data[2]));
 sky130_fd_sc_hd__mux4_2 _399_ (.A0(\memblk.FIFO[0][3] ),
    .A1(\memblk.FIFO[1][3] ),
    .A2(\memblk.FIFO[2][3] ),
    .A3(\memblk.FIFO[3][3] ),
    .S0(_141_),
    .S1(_143_),
    .X(_147_));
 sky130_fd_sc_hd__buf_1 _400_ (.A(_147_),
    .X(F_Data[3]));
 sky130_fd_sc_hd__mux4_2 _401_ (.A0(\memblk.FIFO[0][4] ),
    .A1(\memblk.FIFO[1][4] ),
    .A2(\memblk.FIFO[2][4] ),
    .A3(\memblk.FIFO[3][4] ),
    .S0(_141_),
    .S1(_143_),
    .X(_148_));
 sky130_fd_sc_hd__buf_1 _402_ (.A(_148_),
    .X(F_Data[4]));
 sky130_fd_sc_hd__buf_2 _403_ (.A(_140_),
    .X(_149_));
 sky130_fd_sc_hd__buf_1 _404_ (.A(_142_),
    .X(_150_));
 sky130_fd_sc_hd__mux4_2 _405_ (.A0(\memblk.FIFO[0][5] ),
    .A1(\memblk.FIFO[1][5] ),
    .A2(\memblk.FIFO[2][5] ),
    .A3(\memblk.FIFO[3][5] ),
    .S0(_149_),
    .S1(_150_),
    .X(_151_));
 sky130_fd_sc_hd__buf_1 _406_ (.A(_151_),
    .X(F_Data[5]));
 sky130_fd_sc_hd__mux4_2 _407_ (.A0(\memblk.FIFO[0][6] ),
    .A1(\memblk.FIFO[1][6] ),
    .A2(\memblk.FIFO[2][6] ),
    .A3(\memblk.FIFO[3][6] ),
    .S0(_149_),
    .S1(_150_),
    .X(_152_));
 sky130_fd_sc_hd__buf_1 _408_ (.A(_152_),
    .X(F_Data[6]));
 sky130_fd_sc_hd__mux4_2 _409_ (.A0(\memblk.FIFO[0][7] ),
    .A1(\memblk.FIFO[1][7] ),
    .A2(\memblk.FIFO[2][7] ),
    .A3(\memblk.FIFO[3][7] ),
    .S0(_149_),
    .S1(_150_),
    .X(_153_));
 sky130_fd_sc_hd__buf_1 _410_ (.A(_153_),
    .X(F_Data[7]));
 sky130_fd_sc_hd__mux4_2 _411_ (.A0(\memblk.FIFO[0][8] ),
    .A1(\memblk.FIFO[1][8] ),
    .A2(\memblk.FIFO[2][8] ),
    .A3(\memblk.FIFO[3][8] ),
    .S0(_149_),
    .S1(_150_),
    .X(_154_));
 sky130_fd_sc_hd__buf_1 _412_ (.A(_154_),
    .X(F_Data[8]));
 sky130_fd_sc_hd__mux4_2 _413_ (.A0(\memblk.FIFO[0][9] ),
    .A1(\memblk.FIFO[1][9] ),
    .A2(\memblk.FIFO[2][9] ),
    .A3(\memblk.FIFO[3][9] ),
    .S0(_149_),
    .S1(_150_),
    .X(_155_));
 sky130_fd_sc_hd__buf_1 _414_ (.A(_155_),
    .X(F_Data[9]));
 sky130_fd_sc_hd__mux4_2 _415_ (.A0(\memblk.FIFO[0][10] ),
    .A1(\memblk.FIFO[1][10] ),
    .A2(\memblk.FIFO[2][10] ),
    .A3(\memblk.FIFO[3][10] ),
    .S0(_149_),
    .S1(_150_),
    .X(_156_));
 sky130_fd_sc_hd__buf_1 _416_ (.A(_156_),
    .X(F_Data[10]));
 sky130_fd_sc_hd__buf_1 _417_ (.A(\memblk.rd_addr[0] ),
    .X(_157_));
 sky130_fd_sc_hd__buf_1 _418_ (.A(_142_),
    .X(_158_));
 sky130_fd_sc_hd__mux4_2 _419_ (.A0(\memblk.FIFO[0][11] ),
    .A1(\memblk.FIFO[1][11] ),
    .A2(\memblk.FIFO[2][11] ),
    .A3(\memblk.FIFO[3][11] ),
    .S0(_157_),
    .S1(_158_),
    .X(_159_));
 sky130_fd_sc_hd__buf_1 _420_ (.A(_159_),
    .X(F_Data[11]));
 sky130_fd_sc_hd__mux4_2 _421_ (.A0(\memblk.FIFO[0][12] ),
    .A1(\memblk.FIFO[1][12] ),
    .A2(\memblk.FIFO[2][12] ),
    .A3(\memblk.FIFO[3][12] ),
    .S0(_157_),
    .S1(_158_),
    .X(_160_));
 sky130_fd_sc_hd__buf_1 _422_ (.A(_160_),
    .X(F_Data[12]));
 sky130_fd_sc_hd__mux4_2 _423_ (.A0(\memblk.FIFO[0][13] ),
    .A1(\memblk.FIFO[1][13] ),
    .A2(\memblk.FIFO[2][13] ),
    .A3(\memblk.FIFO[3][13] ),
    .S0(_157_),
    .S1(_158_),
    .X(_161_));
 sky130_fd_sc_hd__buf_1 _424_ (.A(_161_),
    .X(F_Data[13]));
 sky130_fd_sc_hd__mux4_2 _425_ (.A0(\memblk.FIFO[0][14] ),
    .A1(\memblk.FIFO[1][14] ),
    .A2(\memblk.FIFO[2][14] ),
    .A3(\memblk.FIFO[3][14] ),
    .S0(_157_),
    .S1(_158_),
    .X(_162_));
 sky130_fd_sc_hd__buf_1 _426_ (.A(_162_),
    .X(F_Data[14]));
 sky130_fd_sc_hd__mux4_2 _427_ (.A0(\memblk.FIFO[0][15] ),
    .A1(\memblk.FIFO[1][15] ),
    .A2(\memblk.FIFO[2][15] ),
    .A3(\memblk.FIFO[3][15] ),
    .S0(_157_),
    .S1(_158_),
    .X(_163_));
 sky130_fd_sc_hd__buf_1 _428_ (.A(_163_),
    .X(F_Data[15]));
 sky130_fd_sc_hd__mux4_2 _429_ (.A0(\memblk.FIFO[0][16] ),
    .A1(\memblk.FIFO[1][16] ),
    .A2(\memblk.FIFO[2][16] ),
    .A3(\memblk.FIFO[3][16] ),
    .S0(_157_),
    .S1(_158_),
    .X(_164_));
 sky130_fd_sc_hd__buf_1 _430_ (.A(_164_),
    .X(F_Data[16]));
 sky130_fd_sc_hd__buf_2 _431_ (.A(\memblk.rd_addr[0] ),
    .X(_165_));
 sky130_fd_sc_hd__buf_1 _432_ (.A(\memblk.rd_addr[1] ),
    .X(_166_));
 sky130_fd_sc_hd__mux4_2 _433_ (.A0(\memblk.FIFO[0][17] ),
    .A1(\memblk.FIFO[1][17] ),
    .A2(\memblk.FIFO[2][17] ),
    .A3(\memblk.FIFO[3][17] ),
    .S0(_165_),
    .S1(_166_),
    .X(_167_));
 sky130_fd_sc_hd__buf_1 _434_ (.A(_167_),
    .X(F_Data[17]));
 sky130_fd_sc_hd__mux4_2 _435_ (.A0(\memblk.FIFO[0][18] ),
    .A1(\memblk.FIFO[1][18] ),
    .A2(\memblk.FIFO[2][18] ),
    .A3(\memblk.FIFO[3][18] ),
    .S0(_165_),
    .S1(_166_),
    .X(_168_));
 sky130_fd_sc_hd__buf_1 _436_ (.A(_168_),
    .X(F_Data[18]));
 sky130_fd_sc_hd__mux4_2 _437_ (.A0(\memblk.FIFO[0][19] ),
    .A1(\memblk.FIFO[1][19] ),
    .A2(\memblk.FIFO[2][19] ),
    .A3(\memblk.FIFO[3][19] ),
    .S0(_165_),
    .S1(_166_),
    .X(_169_));
 sky130_fd_sc_hd__buf_1 _438_ (.A(_169_),
    .X(F_Data[19]));
 sky130_fd_sc_hd__mux4_2 _439_ (.A0(\memblk.FIFO[0][20] ),
    .A1(\memblk.FIFO[1][20] ),
    .A2(\memblk.FIFO[2][20] ),
    .A3(\memblk.FIFO[3][20] ),
    .S0(_165_),
    .S1(_166_),
    .X(_170_));
 sky130_fd_sc_hd__buf_1 _440_ (.A(_170_),
    .X(F_Data[20]));
 sky130_fd_sc_hd__mux4_2 _441_ (.A0(\memblk.FIFO[0][21] ),
    .A1(\memblk.FIFO[1][21] ),
    .A2(\memblk.FIFO[2][21] ),
    .A3(\memblk.FIFO[3][21] ),
    .S0(_165_),
    .S1(_166_),
    .X(_171_));
 sky130_fd_sc_hd__buf_1 _442_ (.A(_171_),
    .X(F_Data[21]));
 sky130_fd_sc_hd__mux4_2 _443_ (.A0(\memblk.FIFO[0][22] ),
    .A1(\memblk.FIFO[1][22] ),
    .A2(\memblk.FIFO[2][22] ),
    .A3(\memblk.FIFO[3][22] ),
    .S0(_165_),
    .S1(_166_),
    .X(_172_));
 sky130_fd_sc_hd__buf_1 _444_ (.A(_172_),
    .X(F_Data[22]));
 sky130_fd_sc_hd__buf_2 _445_ (.A(\memblk.rd_addr[0] ),
    .X(_173_));
 sky130_fd_sc_hd__buf_1 _446_ (.A(\memblk.rd_addr[1] ),
    .X(_174_));
 sky130_fd_sc_hd__mux4_2 _447_ (.A0(\memblk.FIFO[0][23] ),
    .A1(\memblk.FIFO[1][23] ),
    .A2(\memblk.FIFO[2][23] ),
    .A3(\memblk.FIFO[3][23] ),
    .S0(_173_),
    .S1(_174_),
    .X(_175_));
 sky130_fd_sc_hd__buf_1 _448_ (.A(_175_),
    .X(F_Data[23]));
 sky130_fd_sc_hd__mux4_2 _449_ (.A0(\memblk.FIFO[0][24] ),
    .A1(\memblk.FIFO[1][24] ),
    .A2(\memblk.FIFO[2][24] ),
    .A3(\memblk.FIFO[3][24] ),
    .S0(_173_),
    .S1(_174_),
    .X(_176_));
 sky130_fd_sc_hd__buf_1 _450_ (.A(_176_),
    .X(F_Data[24]));
 sky130_fd_sc_hd__mux4_2 _451_ (.A0(\memblk.FIFO[0][25] ),
    .A1(\memblk.FIFO[1][25] ),
    .A2(\memblk.FIFO[2][25] ),
    .A3(\memblk.FIFO[3][25] ),
    .S0(_173_),
    .S1(_174_),
    .X(_177_));
 sky130_fd_sc_hd__buf_1 _452_ (.A(_177_),
    .X(F_Data[25]));
 sky130_fd_sc_hd__mux4_2 _453_ (.A0(\memblk.FIFO[0][26] ),
    .A1(\memblk.FIFO[1][26] ),
    .A2(\memblk.FIFO[2][26] ),
    .A3(\memblk.FIFO[3][26] ),
    .S0(_173_),
    .S1(_174_),
    .X(_178_));
 sky130_fd_sc_hd__buf_1 _454_ (.A(_178_),
    .X(F_Data[26]));
 sky130_fd_sc_hd__mux4_2 _455_ (.A0(\memblk.FIFO[0][27] ),
    .A1(\memblk.FIFO[1][27] ),
    .A2(\memblk.FIFO[2][27] ),
    .A3(\memblk.FIFO[3][27] ),
    .S0(_173_),
    .S1(_174_),
    .X(_179_));
 sky130_fd_sc_hd__buf_1 _456_ (.A(_179_),
    .X(F_Data[27]));
 sky130_fd_sc_hd__mux4_2 _457_ (.A0(\memblk.FIFO[0][28] ),
    .A1(\memblk.FIFO[1][28] ),
    .A2(\memblk.FIFO[2][28] ),
    .A3(\memblk.FIFO[3][28] ),
    .S0(_173_),
    .S1(_174_),
    .X(_180_));
 sky130_fd_sc_hd__buf_1 _458_ (.A(_180_),
    .X(F_Data[28]));
 sky130_fd_sc_hd__mux4_2 _459_ (.A0(\memblk.FIFO[0][29] ),
    .A1(\memblk.FIFO[1][29] ),
    .A2(\memblk.FIFO[2][29] ),
    .A3(\memblk.FIFO[3][29] ),
    .S0(_140_),
    .S1(_142_),
    .X(_181_));
 sky130_fd_sc_hd__buf_1 _460_ (.A(_181_),
    .X(F_Data[29]));
 sky130_fd_sc_hd__mux4_2 _461_ (.A0(\memblk.FIFO[0][30] ),
    .A1(\memblk.FIFO[1][30] ),
    .A2(\memblk.FIFO[2][30] ),
    .A3(\memblk.FIFO[3][30] ),
    .S0(_140_),
    .S1(_142_),
    .X(_182_));
 sky130_fd_sc_hd__buf_1 _462_ (.A(_182_),
    .X(F_Data[30]));
 sky130_fd_sc_hd__mux4_2 _463_ (.A0(\memblk.FIFO[0][31] ),
    .A1(\memblk.FIFO[1][31] ),
    .A2(\memblk.FIFO[2][31] ),
    .A3(\memblk.FIFO[3][31] ),
    .S0(_140_),
    .S1(_142_),
    .X(_183_));
 sky130_fd_sc_hd__buf_1 _464_ (.A(_183_),
    .X(F_Data[31]));
 sky130_fd_sc_hd__or3b_4 _465_ (.A(FInN),
    .B(\memblk.wr_addr[0] ),
    .C_N(\memblk.wr_addr[1] ),
    .X(_184_));
 sky130_fd_sc_hd__buf_1 _466_ (.A(_184_),
    .X(_185_));
 sky130_fd_sc_hd__buf_2 _467_ (.A(_185_),
    .X(_186_));
 sky130_fd_sc_hd__mux2_2 _468_ (.A0(Data_In[0]),
    .A1(\memblk.FIFO[2][0] ),
    .S(_186_),
    .X(_187_));
 sky130_fd_sc_hd__buf_2 _469_ (.A(_187_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_2 _470_ (.A0(Data_In[1]),
    .A1(\memblk.FIFO[2][1] ),
    .S(_186_),
    .X(_188_));
 sky130_fd_sc_hd__buf_2 _471_ (.A(_188_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_2 _472_ (.A0(Data_In[2]),
    .A1(\memblk.FIFO[2][2] ),
    .S(_186_),
    .X(_189_));
 sky130_fd_sc_hd__buf_2 _473_ (.A(_189_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_2 _474_ (.A0(Data_In[3]),
    .A1(\memblk.FIFO[2][3] ),
    .S(_186_),
    .X(_190_));
 sky130_fd_sc_hd__buf_2 _475_ (.A(_190_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_2 _476_ (.A0(Data_In[4]),
    .A1(\memblk.FIFO[2][4] ),
    .S(_186_),
    .X(_191_));
 sky130_fd_sc_hd__buf_2 _477_ (.A(_191_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_2 _478_ (.A0(Data_In[5]),
    .A1(\memblk.FIFO[2][5] ),
    .S(_186_),
    .X(_192_));
 sky130_fd_sc_hd__buf_2 _479_ (.A(_192_),
    .X(_005_));
 sky130_fd_sc_hd__buf_2 _480_ (.A(_185_),
    .X(_193_));
 sky130_fd_sc_hd__mux2_2 _481_ (.A0(Data_In[6]),
    .A1(\memblk.FIFO[2][6] ),
    .S(_193_),
    .X(_194_));
 sky130_fd_sc_hd__buf_2 _482_ (.A(_194_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_2 _483_ (.A0(Data_In[7]),
    .A1(\memblk.FIFO[2][7] ),
    .S(_193_),
    .X(_195_));
 sky130_fd_sc_hd__buf_2 _484_ (.A(_195_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_2 _485_ (.A0(Data_In[8]),
    .A1(\memblk.FIFO[2][8] ),
    .S(_193_),
    .X(_196_));
 sky130_fd_sc_hd__buf_2 _486_ (.A(_196_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_2 _487_ (.A0(Data_In[9]),
    .A1(\memblk.FIFO[2][9] ),
    .S(_193_),
    .X(_197_));
 sky130_fd_sc_hd__buf_2 _488_ (.A(_197_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_2 _489_ (.A0(Data_In[10]),
    .A1(\memblk.FIFO[2][10] ),
    .S(_193_),
    .X(_198_));
 sky130_fd_sc_hd__buf_2 _490_ (.A(_198_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_2 _491_ (.A0(Data_In[11]),
    .A1(\memblk.FIFO[2][11] ),
    .S(_193_),
    .X(_199_));
 sky130_fd_sc_hd__buf_2 _492_ (.A(_199_),
    .X(_011_));
 sky130_fd_sc_hd__buf_2 _493_ (.A(_185_),
    .X(_200_));
 sky130_fd_sc_hd__mux2_2 _494_ (.A0(Data_In[12]),
    .A1(\memblk.FIFO[2][12] ),
    .S(_200_),
    .X(_201_));
 sky130_fd_sc_hd__buf_2 _495_ (.A(_201_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_2 _496_ (.A0(Data_In[13]),
    .A1(\memblk.FIFO[2][13] ),
    .S(_200_),
    .X(_202_));
 sky130_fd_sc_hd__buf_2 _497_ (.A(_202_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_2 _498_ (.A0(Data_In[14]),
    .A1(\memblk.FIFO[2][14] ),
    .S(_200_),
    .X(_203_));
 sky130_fd_sc_hd__buf_2 _499_ (.A(_203_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_2 _500_ (.A0(Data_In[15]),
    .A1(\memblk.FIFO[2][15] ),
    .S(_200_),
    .X(_204_));
 sky130_fd_sc_hd__buf_2 _501_ (.A(_204_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_2 _502_ (.A0(Data_In[16]),
    .A1(\memblk.FIFO[2][16] ),
    .S(_200_),
    .X(_205_));
 sky130_fd_sc_hd__buf_2 _503_ (.A(_205_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_2 _504_ (.A0(Data_In[17]),
    .A1(\memblk.FIFO[2][17] ),
    .S(_200_),
    .X(_206_));
 sky130_fd_sc_hd__buf_2 _505_ (.A(_206_),
    .X(_017_));
 sky130_fd_sc_hd__buf_2 _506_ (.A(_185_),
    .X(_207_));
 sky130_fd_sc_hd__mux2_2 _507_ (.A0(Data_In[18]),
    .A1(\memblk.FIFO[2][18] ),
    .S(_207_),
    .X(_208_));
 sky130_fd_sc_hd__buf_2 _508_ (.A(_208_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_2 _509_ (.A0(Data_In[19]),
    .A1(\memblk.FIFO[2][19] ),
    .S(_207_),
    .X(_209_));
 sky130_fd_sc_hd__buf_2 _510_ (.A(_209_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_2 _511_ (.A0(Data_In[20]),
    .A1(\memblk.FIFO[2][20] ),
    .S(_207_),
    .X(_210_));
 sky130_fd_sc_hd__buf_2 _512_ (.A(_210_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_2 _513_ (.A0(Data_In[21]),
    .A1(\memblk.FIFO[2][21] ),
    .S(_207_),
    .X(_211_));
 sky130_fd_sc_hd__buf_2 _514_ (.A(_211_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_2 _515_ (.A0(Data_In[22]),
    .A1(\memblk.FIFO[2][22] ),
    .S(_207_),
    .X(_212_));
 sky130_fd_sc_hd__buf_2 _516_ (.A(_212_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_2 _517_ (.A0(Data_In[23]),
    .A1(\memblk.FIFO[2][23] ),
    .S(_207_),
    .X(_213_));
 sky130_fd_sc_hd__buf_2 _518_ (.A(_213_),
    .X(_023_));
 sky130_fd_sc_hd__buf_1 _519_ (.A(_184_),
    .X(_214_));
 sky130_fd_sc_hd__mux2_2 _520_ (.A0(Data_In[24]),
    .A1(\memblk.FIFO[2][24] ),
    .S(_214_),
    .X(_215_));
 sky130_fd_sc_hd__buf_1 _521_ (.A(_215_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_2 _522_ (.A0(Data_In[25]),
    .A1(\memblk.FIFO[2][25] ),
    .S(_214_),
    .X(_216_));
 sky130_fd_sc_hd__buf_1 _523_ (.A(_216_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_2 _524_ (.A0(Data_In[26]),
    .A1(\memblk.FIFO[2][26] ),
    .S(_214_),
    .X(_217_));
 sky130_fd_sc_hd__buf_1 _525_ (.A(_217_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_2 _526_ (.A0(Data_In[27]),
    .A1(\memblk.FIFO[2][27] ),
    .S(_214_),
    .X(_218_));
 sky130_fd_sc_hd__buf_1 _527_ (.A(_218_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_2 _528_ (.A0(Data_In[28]),
    .A1(\memblk.FIFO[2][28] ),
    .S(_214_),
    .X(_219_));
 sky130_fd_sc_hd__buf_1 _529_ (.A(_219_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_2 _530_ (.A0(Data_In[29]),
    .A1(\memblk.FIFO[2][29] ),
    .S(_214_),
    .X(_220_));
 sky130_fd_sc_hd__buf_1 _531_ (.A(_220_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_2 _532_ (.A0(Data_In[30]),
    .A1(\memblk.FIFO[2][30] ),
    .S(_185_),
    .X(_221_));
 sky130_fd_sc_hd__buf_1 _533_ (.A(_221_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_2 _534_ (.A0(Data_In[31]),
    .A1(\memblk.FIFO[2][31] ),
    .S(_185_),
    .X(_222_));
 sky130_fd_sc_hd__buf_1 _535_ (.A(_222_),
    .X(_031_));
 sky130_fd_sc_hd__buf_1 _536_ (.A(FClrN),
    .X(_223_));
 sky130_fd_sc_hd__nand2b_2 _537_ (.A_N(FInN),
    .B(\memblk.wr_addr[0] ),
    .Y(_224_));
 sky130_fd_sc_hd__bufinv_8 _538_ (.A(FInN),
    .Y(_225_));
 sky130_fd_sc_hd__or2_2 _539_ (.A(_225_),
    .B(\memblk.wr_addr[0] ),
    .X(_226_));
 sky130_fd_sc_hd__and3_2 _540_ (.A(_223_),
    .B(_224_),
    .C(_226_),
    .X(_227_));
 sky130_fd_sc_hd__buf_1 _541_ (.A(_227_),
    .X(_032_));
 sky130_fd_sc_hd__or2_4 _542_ (.A(\memblk.wr_addr[1] ),
    .B(_224_),
    .X(_228_));
 sky130_fd_sc_hd__buf_1 _543_ (.A(_228_),
    .X(_229_));
 sky130_fd_sc_hd__buf_2 _544_ (.A(_229_),
    .X(_230_));
 sky130_fd_sc_hd__nand2_2 _545_ (.A(\memblk.wr_addr[1] ),
    .B(_224_),
    .Y(_231_));
 sky130_fd_sc_hd__inv_2 _546_ (.A(_223_),
    .Y(_232_));
 sky130_fd_sc_hd__a21oi_2 _547_ (.A1(_230_),
    .A2(_231_),
    .B1(_232_),
    .Y(_033_));
 sky130_fd_sc_hd__or3_4 _548_ (.A(FInN),
    .B(\memblk.wr_addr[0] ),
    .C(\memblk.wr_addr[1] ),
    .X(_233_));
 sky130_fd_sc_hd__buf_1 _549_ (.A(_233_),
    .X(_234_));
 sky130_fd_sc_hd__buf_2 _550_ (.A(_234_),
    .X(_235_));
 sky130_fd_sc_hd__mux2_2 _551_ (.A0(Data_In[0]),
    .A1(\memblk.FIFO[0][0] ),
    .S(_235_),
    .X(_236_));
 sky130_fd_sc_hd__buf_1 _552_ (.A(_236_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_2 _553_ (.A0(Data_In[1]),
    .A1(\memblk.FIFO[0][1] ),
    .S(_235_),
    .X(_237_));
 sky130_fd_sc_hd__buf_1 _554_ (.A(_237_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_2 _555_ (.A0(Data_In[2]),
    .A1(\memblk.FIFO[0][2] ),
    .S(_235_),
    .X(_238_));
 sky130_fd_sc_hd__buf_1 _556_ (.A(_238_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_2 _557_ (.A0(Data_In[3]),
    .A1(\memblk.FIFO[0][3] ),
    .S(_235_),
    .X(_239_));
 sky130_fd_sc_hd__buf_1 _558_ (.A(_239_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_2 _559_ (.A0(Data_In[4]),
    .A1(\memblk.FIFO[0][4] ),
    .S(_235_),
    .X(_240_));
 sky130_fd_sc_hd__buf_1 _560_ (.A(_240_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_2 _561_ (.A0(Data_In[5]),
    .A1(\memblk.FIFO[0][5] ),
    .S(_235_),
    .X(_241_));
 sky130_fd_sc_hd__buf_1 _562_ (.A(_241_),
    .X(_039_));
 sky130_fd_sc_hd__buf_1 _563_ (.A(_234_),
    .X(_242_));
 sky130_fd_sc_hd__mux2_2 _564_ (.A0(Data_In[6]),
    .A1(\memblk.FIFO[0][6] ),
    .S(_242_),
    .X(_243_));
 sky130_fd_sc_hd__buf_2 _565_ (.A(_243_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_2 _566_ (.A0(Data_In[7]),
    .A1(\memblk.FIFO[0][7] ),
    .S(_242_),
    .X(_244_));
 sky130_fd_sc_hd__buf_2 _567_ (.A(_244_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_2 _568_ (.A0(Data_In[8]),
    .A1(\memblk.FIFO[0][8] ),
    .S(_242_),
    .X(_245_));
 sky130_fd_sc_hd__buf_2 _569_ (.A(_245_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_2 _570_ (.A0(Data_In[9]),
    .A1(\memblk.FIFO[0][9] ),
    .S(_242_),
    .X(_246_));
 sky130_fd_sc_hd__buf_2 _571_ (.A(_246_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_2 _572_ (.A0(Data_In[10]),
    .A1(\memblk.FIFO[0][10] ),
    .S(_242_),
    .X(_247_));
 sky130_fd_sc_hd__buf_2 _573_ (.A(_247_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_2 _574_ (.A0(Data_In[11]),
    .A1(\memblk.FIFO[0][11] ),
    .S(_242_),
    .X(_248_));
 sky130_fd_sc_hd__buf_2 _575_ (.A(_248_),
    .X(_045_));
 sky130_fd_sc_hd__buf_2 _576_ (.A(_234_),
    .X(_249_));
 sky130_fd_sc_hd__mux2_2 _577_ (.A0(Data_In[12]),
    .A1(\memblk.FIFO[0][12] ),
    .S(_249_),
    .X(_250_));
 sky130_fd_sc_hd__buf_1 _578_ (.A(_250_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_2 _579_ (.A0(Data_In[13]),
    .A1(\memblk.FIFO[0][13] ),
    .S(_249_),
    .X(_251_));
 sky130_fd_sc_hd__buf_1 _580_ (.A(_251_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_2 _581_ (.A0(Data_In[14]),
    .A1(\memblk.FIFO[0][14] ),
    .S(_249_),
    .X(_252_));
 sky130_fd_sc_hd__buf_1 _582_ (.A(_252_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_2 _583_ (.A0(Data_In[15]),
    .A1(\memblk.FIFO[0][15] ),
    .S(_249_),
    .X(_253_));
 sky130_fd_sc_hd__buf_1 _584_ (.A(_253_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_2 _585_ (.A0(Data_In[16]),
    .A1(\memblk.FIFO[0][16] ),
    .S(_249_),
    .X(_254_));
 sky130_fd_sc_hd__buf_1 _586_ (.A(_254_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_2 _587_ (.A0(Data_In[17]),
    .A1(\memblk.FIFO[0][17] ),
    .S(_249_),
    .X(_255_));
 sky130_fd_sc_hd__buf_1 _588_ (.A(_255_),
    .X(_051_));
 sky130_fd_sc_hd__buf_2 _589_ (.A(_234_),
    .X(_256_));
 sky130_fd_sc_hd__mux2_2 _590_ (.A0(Data_In[18]),
    .A1(\memblk.FIFO[0][18] ),
    .S(_256_),
    .X(_257_));
 sky130_fd_sc_hd__buf_1 _591_ (.A(_257_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_2 _592_ (.A0(Data_In[19]),
    .A1(\memblk.FIFO[0][19] ),
    .S(_256_),
    .X(_258_));
 sky130_fd_sc_hd__buf_1 _593_ (.A(_258_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_2 _594_ (.A0(Data_In[20]),
    .A1(\memblk.FIFO[0][20] ),
    .S(_256_),
    .X(_259_));
 sky130_fd_sc_hd__buf_1 _595_ (.A(_259_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_2 _596_ (.A0(Data_In[21]),
    .A1(\memblk.FIFO[0][21] ),
    .S(_256_),
    .X(_260_));
 sky130_fd_sc_hd__buf_1 _597_ (.A(_260_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_2 _598_ (.A0(Data_In[22]),
    .A1(\memblk.FIFO[0][22] ),
    .S(_256_),
    .X(_261_));
 sky130_fd_sc_hd__buf_1 _599_ (.A(_261_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_2 _600_ (.A0(Data_In[23]),
    .A1(\memblk.FIFO[0][23] ),
    .S(_256_),
    .X(_262_));
 sky130_fd_sc_hd__buf_1 _601_ (.A(_262_),
    .X(_057_));
 sky130_fd_sc_hd__buf_1 _602_ (.A(_233_),
    .X(_263_));
 sky130_fd_sc_hd__mux2_2 _603_ (.A0(Data_In[24]),
    .A1(\memblk.FIFO[0][24] ),
    .S(_263_),
    .X(_264_));
 sky130_fd_sc_hd__buf_1 _604_ (.A(_264_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_2 _605_ (.A0(Data_In[25]),
    .A1(\memblk.FIFO[0][25] ),
    .S(_263_),
    .X(_265_));
 sky130_fd_sc_hd__buf_1 _606_ (.A(_265_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_2 _607_ (.A0(Data_In[26]),
    .A1(\memblk.FIFO[0][26] ),
    .S(_263_),
    .X(_266_));
 sky130_fd_sc_hd__buf_1 _608_ (.A(_266_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_2 _609_ (.A0(Data_In[27]),
    .A1(\memblk.FIFO[0][27] ),
    .S(_263_),
    .X(_267_));
 sky130_fd_sc_hd__buf_1 _610_ (.A(_267_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_2 _611_ (.A0(Data_In[28]),
    .A1(\memblk.FIFO[0][28] ),
    .S(_263_),
    .X(_268_));
 sky130_fd_sc_hd__buf_1 _612_ (.A(_268_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_2 _613_ (.A0(Data_In[29]),
    .A1(\memblk.FIFO[0][29] ),
    .S(_263_),
    .X(_269_));
 sky130_fd_sc_hd__buf_1 _614_ (.A(_269_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_2 _615_ (.A0(Data_In[30]),
    .A1(\memblk.FIFO[0][30] ),
    .S(_234_),
    .X(_270_));
 sky130_fd_sc_hd__buf_1 _616_ (.A(_270_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_2 _617_ (.A0(Data_In[31]),
    .A1(\memblk.FIFO[0][31] ),
    .S(_234_),
    .X(_271_));
 sky130_fd_sc_hd__buf_1 _618_ (.A(_271_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_2 _619_ (.A0(Data_In[0]),
    .A1(\memblk.FIFO[1][0] ),
    .S(_230_),
    .X(_272_));
 sky130_fd_sc_hd__buf_2 _620_ (.A(_272_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_2 _621_ (.A0(Data_In[1]),
    .A1(\memblk.FIFO[1][1] ),
    .S(_230_),
    .X(_273_));
 sky130_fd_sc_hd__buf_2 _622_ (.A(_273_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_2 _623_ (.A0(Data_In[2]),
    .A1(\memblk.FIFO[1][2] ),
    .S(_230_),
    .X(_274_));
 sky130_fd_sc_hd__buf_2 _624_ (.A(_274_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_2 _625_ (.A0(Data_In[3]),
    .A1(\memblk.FIFO[1][3] ),
    .S(_230_),
    .X(_275_));
 sky130_fd_sc_hd__buf_2 _626_ (.A(_275_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_2 _627_ (.A0(Data_In[4]),
    .A1(\memblk.FIFO[1][4] ),
    .S(_230_),
    .X(_276_));
 sky130_fd_sc_hd__buf_2 _628_ (.A(_276_),
    .X(_070_));
 sky130_fd_sc_hd__buf_2 _629_ (.A(_229_),
    .X(_277_));
 sky130_fd_sc_hd__mux2_2 _630_ (.A0(Data_In[5]),
    .A1(\memblk.FIFO[1][5] ),
    .S(_277_),
    .X(_278_));
 sky130_fd_sc_hd__buf_2 _631_ (.A(_278_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_2 _632_ (.A0(Data_In[6]),
    .A1(\memblk.FIFO[1][6] ),
    .S(_277_),
    .X(_279_));
 sky130_fd_sc_hd__buf_2 _633_ (.A(_279_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_2 _634_ (.A0(Data_In[7]),
    .A1(\memblk.FIFO[1][7] ),
    .S(_277_),
    .X(_280_));
 sky130_fd_sc_hd__buf_2 _635_ (.A(_280_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_2 _636_ (.A0(Data_In[8]),
    .A1(\memblk.FIFO[1][8] ),
    .S(_277_),
    .X(_281_));
 sky130_fd_sc_hd__buf_2 _637_ (.A(_281_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_2 _638_ (.A0(Data_In[9]),
    .A1(\memblk.FIFO[1][9] ),
    .S(_277_),
    .X(_282_));
 sky130_fd_sc_hd__buf_2 _639_ (.A(_282_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_2 _640_ (.A0(Data_In[10]),
    .A1(\memblk.FIFO[1][10] ),
    .S(_277_),
    .X(_283_));
 sky130_fd_sc_hd__buf_2 _641_ (.A(_283_),
    .X(_076_));
 sky130_fd_sc_hd__buf_2 _642_ (.A(_229_),
    .X(_284_));
 sky130_fd_sc_hd__mux2_2 _643_ (.A0(Data_In[11]),
    .A1(\memblk.FIFO[1][11] ),
    .S(_284_),
    .X(_285_));
 sky130_fd_sc_hd__buf_2 _644_ (.A(_285_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_2 _645_ (.A0(Data_In[12]),
    .A1(\memblk.FIFO[1][12] ),
    .S(_284_),
    .X(_286_));
 sky130_fd_sc_hd__buf_2 _646_ (.A(_286_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_2 _647_ (.A0(Data_In[13]),
    .A1(\memblk.FIFO[1][13] ),
    .S(_284_),
    .X(_287_));
 sky130_fd_sc_hd__buf_2 _648_ (.A(_287_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_2 _649_ (.A0(Data_In[14]),
    .A1(\memblk.FIFO[1][14] ),
    .S(_284_),
    .X(_288_));
 sky130_fd_sc_hd__buf_2 _650_ (.A(_288_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_2 _651_ (.A0(Data_In[15]),
    .A1(\memblk.FIFO[1][15] ),
    .S(_284_),
    .X(_289_));
 sky130_fd_sc_hd__buf_2 _652_ (.A(_289_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_2 _653_ (.A0(Data_In[16]),
    .A1(\memblk.FIFO[1][16] ),
    .S(_284_),
    .X(_290_));
 sky130_fd_sc_hd__buf_2 _654_ (.A(_290_),
    .X(_082_));
 sky130_fd_sc_hd__buf_1 _655_ (.A(_228_),
    .X(_291_));
 sky130_fd_sc_hd__mux2_2 _656_ (.A0(Data_In[17]),
    .A1(\memblk.FIFO[1][17] ),
    .S(_291_),
    .X(_292_));
 sky130_fd_sc_hd__buf_1 _657_ (.A(_292_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_2 _658_ (.A0(Data_In[18]),
    .A1(\memblk.FIFO[1][18] ),
    .S(_291_),
    .X(_293_));
 sky130_fd_sc_hd__buf_1 _659_ (.A(_293_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_2 _660_ (.A0(Data_In[19]),
    .A1(\memblk.FIFO[1][19] ),
    .S(_291_),
    .X(_294_));
 sky130_fd_sc_hd__buf_1 _661_ (.A(_294_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_2 _662_ (.A0(Data_In[20]),
    .A1(\memblk.FIFO[1][20] ),
    .S(_291_),
    .X(_295_));
 sky130_fd_sc_hd__buf_1 _663_ (.A(_295_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_2 _664_ (.A0(Data_In[21]),
    .A1(\memblk.FIFO[1][21] ),
    .S(_291_),
    .X(_296_));
 sky130_fd_sc_hd__buf_1 _665_ (.A(_296_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_2 _666_ (.A0(Data_In[22]),
    .A1(\memblk.FIFO[1][22] ),
    .S(_291_),
    .X(_297_));
 sky130_fd_sc_hd__buf_1 _667_ (.A(_297_),
    .X(_088_));
 sky130_fd_sc_hd__buf_1 _668_ (.A(_228_),
    .X(_298_));
 sky130_fd_sc_hd__mux2_2 _669_ (.A0(Data_In[23]),
    .A1(\memblk.FIFO[1][23] ),
    .S(_298_),
    .X(_299_));
 sky130_fd_sc_hd__buf_1 _670_ (.A(_299_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_2 _671_ (.A0(Data_In[24]),
    .A1(\memblk.FIFO[1][24] ),
    .S(_298_),
    .X(_300_));
 sky130_fd_sc_hd__buf_1 _672_ (.A(_300_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_2 _673_ (.A0(Data_In[25]),
    .A1(\memblk.FIFO[1][25] ),
    .S(_298_),
    .X(_301_));
 sky130_fd_sc_hd__buf_1 _674_ (.A(_301_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_2 _675_ (.A0(Data_In[26]),
    .A1(\memblk.FIFO[1][26] ),
    .S(_298_),
    .X(_302_));
 sky130_fd_sc_hd__buf_1 _676_ (.A(_302_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_2 _677_ (.A0(Data_In[27]),
    .A1(\memblk.FIFO[1][27] ),
    .S(_298_),
    .X(_303_));
 sky130_fd_sc_hd__buf_1 _678_ (.A(_303_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_2 _679_ (.A0(Data_In[28]),
    .A1(\memblk.FIFO[1][28] ),
    .S(_298_),
    .X(_304_));
 sky130_fd_sc_hd__buf_1 _680_ (.A(_304_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_2 _681_ (.A0(Data_In[29]),
    .A1(\memblk.FIFO[1][29] ),
    .S(_229_),
    .X(_305_));
 sky130_fd_sc_hd__buf_1 _682_ (.A(_305_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_2 _683_ (.A0(Data_In[30]),
    .A1(\memblk.FIFO[1][30] ),
    .S(_229_),
    .X(_306_));
 sky130_fd_sc_hd__buf_1 _684_ (.A(_306_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_2 _685_ (.A0(Data_In[31]),
    .A1(\memblk.FIFO[1][31] ),
    .S(_229_),
    .X(_307_));
 sky130_fd_sc_hd__buf_1 _686_ (.A(_307_),
    .X(_097_));
 sky130_fd_sc_hd__and3_2 _687_ (.A(_225_),
    .B(\memblk.wr_addr[0] ),
    .C(\memblk.wr_addr[1] ),
    .X(_308_));
 sky130_fd_sc_hd__buf_1 _688_ (.A(_308_),
    .X(_309_));
 sky130_fd_sc_hd__buf_2 _689_ (.A(_309_),
    .X(_310_));
 sky130_fd_sc_hd__mux2_2 _690_ (.A0(\memblk.FIFO[3][0] ),
    .A1(Data_In[0]),
    .S(_310_),
    .X(_311_));
 sky130_fd_sc_hd__buf_2 _691_ (.A(_311_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_2 _692_ (.A0(\memblk.FIFO[3][1] ),
    .A1(Data_In[1]),
    .S(_310_),
    .X(_312_));
 sky130_fd_sc_hd__buf_2 _693_ (.A(_312_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_2 _694_ (.A0(\memblk.FIFO[3][2] ),
    .A1(Data_In[2]),
    .S(_310_),
    .X(_313_));
 sky130_fd_sc_hd__buf_2 _695_ (.A(_313_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_2 _696_ (.A0(\memblk.FIFO[3][3] ),
    .A1(Data_In[3]),
    .S(_310_),
    .X(_314_));
 sky130_fd_sc_hd__buf_2 _697_ (.A(_314_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_2 _698_ (.A0(\memblk.FIFO[3][4] ),
    .A1(Data_In[4]),
    .S(_310_),
    .X(_315_));
 sky130_fd_sc_hd__buf_2 _699_ (.A(_315_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_2 _700_ (.A0(\memblk.FIFO[3][5] ),
    .A1(Data_In[5]),
    .S(_310_),
    .X(_316_));
 sky130_fd_sc_hd__buf_2 _701_ (.A(_316_),
    .X(_103_));
 sky130_fd_sc_hd__buf_2 _702_ (.A(_309_),
    .X(_317_));
 sky130_fd_sc_hd__mux2_2 _703_ (.A0(\memblk.FIFO[3][6] ),
    .A1(Data_In[6]),
    .S(_317_),
    .X(_318_));
 sky130_fd_sc_hd__buf_2 _704_ (.A(_318_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_2 _705_ (.A0(\memblk.FIFO[3][7] ),
    .A1(Data_In[7]),
    .S(_317_),
    .X(_319_));
 sky130_fd_sc_hd__buf_2 _706_ (.A(_319_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_2 _707_ (.A0(\memblk.FIFO[3][8] ),
    .A1(Data_In[8]),
    .S(_317_),
    .X(_320_));
 sky130_fd_sc_hd__buf_2 _708_ (.A(_320_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_2 _709_ (.A0(\memblk.FIFO[3][9] ),
    .A1(Data_In[9]),
    .S(_317_),
    .X(_321_));
 sky130_fd_sc_hd__buf_2 _710_ (.A(_321_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_2 _711_ (.A0(\memblk.FIFO[3][10] ),
    .A1(Data_In[10]),
    .S(_317_),
    .X(_322_));
 sky130_fd_sc_hd__buf_2 _712_ (.A(_322_),
    .X(_108_));
 sky130_fd_sc_hd__mux2_2 _713_ (.A0(\memblk.FIFO[3][11] ),
    .A1(Data_In[11]),
    .S(_317_),
    .X(_323_));
 sky130_fd_sc_hd__buf_2 _714_ (.A(_323_),
    .X(_109_));
 sky130_fd_sc_hd__buf_2 _715_ (.A(_309_),
    .X(_324_));
 sky130_fd_sc_hd__mux2_2 _716_ (.A0(\memblk.FIFO[3][12] ),
    .A1(Data_In[12]),
    .S(_324_),
    .X(_325_));
 sky130_fd_sc_hd__buf_2 _717_ (.A(_325_),
    .X(_110_));
 sky130_fd_sc_hd__mux2_2 _718_ (.A0(\memblk.FIFO[3][13] ),
    .A1(Data_In[13]),
    .S(_324_),
    .X(_326_));
 sky130_fd_sc_hd__buf_2 _719_ (.A(_326_),
    .X(_111_));
 sky130_fd_sc_hd__mux2_2 _720_ (.A0(\memblk.FIFO[3][14] ),
    .A1(Data_In[14]),
    .S(_324_),
    .X(_327_));
 sky130_fd_sc_hd__buf_2 _721_ (.A(_327_),
    .X(_112_));
 sky130_fd_sc_hd__mux2_2 _722_ (.A0(\memblk.FIFO[3][15] ),
    .A1(Data_In[15]),
    .S(_324_),
    .X(_328_));
 sky130_fd_sc_hd__buf_2 _723_ (.A(_328_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_2 _724_ (.A0(\memblk.FIFO[3][16] ),
    .A1(Data_In[16]),
    .S(_324_),
    .X(_329_));
 sky130_fd_sc_hd__buf_2 _725_ (.A(_329_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_2 _726_ (.A0(\memblk.FIFO[3][17] ),
    .A1(Data_In[17]),
    .S(_324_),
    .X(_330_));
 sky130_fd_sc_hd__buf_2 _727_ (.A(_330_),
    .X(_115_));
 sky130_fd_sc_hd__buf_2 _728_ (.A(_309_),
    .X(_331_));
 sky130_fd_sc_hd__mux2_2 _729_ (.A0(\memblk.FIFO[3][18] ),
    .A1(Data_In[18]),
    .S(_331_),
    .X(_332_));
 sky130_fd_sc_hd__buf_2 _730_ (.A(_332_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_2 _731_ (.A0(\memblk.FIFO[3][19] ),
    .A1(Data_In[19]),
    .S(_331_),
    .X(_333_));
 sky130_fd_sc_hd__buf_2 _732_ (.A(_333_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_2 _733_ (.A0(\memblk.FIFO[3][20] ),
    .A1(Data_In[20]),
    .S(_331_),
    .X(_334_));
 sky130_fd_sc_hd__buf_2 _734_ (.A(_334_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_2 _735_ (.A0(\memblk.FIFO[3][21] ),
    .A1(Data_In[21]),
    .S(_331_),
    .X(_335_));
 sky130_fd_sc_hd__buf_2 _736_ (.A(_335_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_2 _737_ (.A0(\memblk.FIFO[3][22] ),
    .A1(Data_In[22]),
    .S(_331_),
    .X(_336_));
 sky130_fd_sc_hd__buf_2 _738_ (.A(_336_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_2 _739_ (.A0(\memblk.FIFO[3][23] ),
    .A1(Data_In[23]),
    .S(_331_),
    .X(_337_));
 sky130_fd_sc_hd__buf_2 _740_ (.A(_337_),
    .X(_121_));
 sky130_fd_sc_hd__buf_2 _741_ (.A(_308_),
    .X(_338_));
 sky130_fd_sc_hd__mux2_2 _742_ (.A0(\memblk.FIFO[3][24] ),
    .A1(Data_In[24]),
    .S(_338_),
    .X(_339_));
 sky130_fd_sc_hd__buf_1 _743_ (.A(_339_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_2 _744_ (.A0(\memblk.FIFO[3][25] ),
    .A1(Data_In[25]),
    .S(_338_),
    .X(_340_));
 sky130_fd_sc_hd__buf_1 _745_ (.A(_340_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_2 _746_ (.A0(\memblk.FIFO[3][26] ),
    .A1(Data_In[26]),
    .S(_338_),
    .X(_341_));
 sky130_fd_sc_hd__buf_1 _747_ (.A(_341_),
    .X(_124_));
 sky130_fd_sc_hd__mux2_2 _748_ (.A0(\memblk.FIFO[3][27] ),
    .A1(Data_In[27]),
    .S(_338_),
    .X(_342_));
 sky130_fd_sc_hd__buf_1 _749_ (.A(_342_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_2 _750_ (.A0(\memblk.FIFO[3][28] ),
    .A1(Data_In[28]),
    .S(_338_),
    .X(_343_));
 sky130_fd_sc_hd__buf_1 _751_ (.A(_343_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_2 _752_ (.A0(\memblk.FIFO[3][29] ),
    .A1(Data_In[29]),
    .S(_338_),
    .X(_344_));
 sky130_fd_sc_hd__buf_1 _753_ (.A(_344_),
    .X(_127_));
 sky130_fd_sc_hd__mux2_2 _754_ (.A0(\memblk.FIFO[3][30] ),
    .A1(Data_In[30]),
    .S(_309_),
    .X(_345_));
 sky130_fd_sc_hd__buf_1 _755_ (.A(_345_),
    .X(_128_));
 sky130_fd_sc_hd__mux2_2 _756_ (.A0(\memblk.FIFO[3][31] ),
    .A1(Data_In[31]),
    .S(_309_),
    .X(_346_));
 sky130_fd_sc_hd__buf_1 _757_ (.A(_346_),
    .X(_129_));
 sky130_fd_sc_hd__inv_2 _758_ (.A(FOutN),
    .Y(_347_));
 sky130_fd_sc_hd__buf_6 _759_ (.A(FInN),
    .X(_348_));
 sky130_fd_sc_hd__buf_1 _760_ (.A(_348_),
    .X(_349_));
 sky130_fd_sc_hd__o21ai_2 _761_ (.A1(F_LastN),
    .A2(_349_),
    .B1(F_FullN),
    .Y(_350_));
 sky130_fd_sc_hd__or3b_2 _762_ (.A(_347_),
    .B(_232_),
    .C_N(_350_),
    .X(_351_));
 sky130_fd_sc_hd__buf_1 _763_ (.A(_351_),
    .X(_130_));
 sky130_fd_sc_hd__buf_1 _764_ (.A(FOutN),
    .X(_352_));
 sky130_fd_sc_hd__nor2_2 _765_ (.A(_352_),
    .B(_350_),
    .Y(_353_));
 sky130_fd_sc_hd__buf_2 _766_ (.A(\fcounter[0] ),
    .X(_354_));
 sky130_fd_sc_hd__or4b_4 _767_ (.A(_348_),
    .B(_354_),
    .C(\fcounter[2] ),
    .D_N(\fcounter[1] ),
    .X(_355_));
 sky130_fd_sc_hd__o211a_2 _768_ (.A1(F_LastN),
    .A2(_225_),
    .B1(_355_),
    .C1(_352_),
    .X(_356_));
 sky130_fd_sc_hd__or3_4 _769_ (.A(_232_),
    .B(_353_),
    .C(_356_),
    .X(_357_));
 sky130_fd_sc_hd__buf_2 _770_ (.A(_357_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_2 _771_ (.A0(F_SLastN),
    .A1(F_LastN),
    .S(_349_),
    .X(_358_));
 sky130_fd_sc_hd__buf_1 _772_ (.A(\fcounter[2] ),
    .X(_359_));
 sky130_fd_sc_hd__or4b_2 _773_ (.A(_348_),
    .B(\fcounter[1] ),
    .C(_359_),
    .D_N(_354_),
    .X(_360_));
 sky130_fd_sc_hd__o211a_2 _774_ (.A1(_225_),
    .A2(F_SLastN),
    .B1(_360_),
    .C1(_352_),
    .X(_361_));
 sky130_fd_sc_hd__a211o_4 _775_ (.A1(_347_),
    .A2(_358_),
    .B1(_361_),
    .C1(_232_),
    .X(_132_));
 sky130_fd_sc_hd__inv_2 _776_ (.A(F_FirstN),
    .Y(_362_));
 sky130_fd_sc_hd__nor2_2 _777_ (.A(_349_),
    .B(F_EmptyN),
    .Y(_363_));
 sky130_fd_sc_hd__a31o_2 _778_ (.A1(_352_),
    .A2(_349_),
    .A3(_362_),
    .B1(_363_),
    .X(_364_));
 sky130_fd_sc_hd__nand4bb_2 _779_ (.A_N(_354_),
    .B_N(_359_),
    .C(_349_),
    .D(\fcounter[1] ),
    .Y(_365_));
 sky130_fd_sc_hd__or2_2 _780_ (.A(_349_),
    .B(F_FirstN),
    .X(_366_));
 sky130_fd_sc_hd__a21oi_2 _781_ (.A1(_365_),
    .A2(_366_),
    .B1(_352_),
    .Y(_367_));
 sky130_fd_sc_hd__o21ai_2 _782_ (.A1(_364_),
    .A2(_367_),
    .B1(_223_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2_2 _783_ (.A0(F_EmptyN),
    .A1(_363_),
    .S(_223_),
    .X(_368_));
 sky130_fd_sc_hd__buf_1 _784_ (.A(_368_),
    .X(_134_));
 sky130_fd_sc_hd__and2_2 _785_ (.A(_223_),
    .B(_354_),
    .X(_369_));
 sky130_fd_sc_hd__nor2_2 _786_ (.A(_232_),
    .B(_354_),
    .Y(_370_));
 sky130_fd_sc_hd__and3b_2 _787_ (.A_N(FOutN),
    .B(_348_),
    .C(F_EmptyN),
    .X(_371_));
 sky130_fd_sc_hd__a31o_2 _788_ (.A1(F_FullN),
    .A2(FOutN),
    .A3(_225_),
    .B1(_371_),
    .X(_372_));
 sky130_fd_sc_hd__mux2_2 _789_ (.A0(_369_),
    .A1(_370_),
    .S(_372_),
    .X(_373_));
 sky130_fd_sc_hd__buf_1 _790_ (.A(_373_),
    .X(_135_));
 sky130_fd_sc_hd__and2b_2 _791_ (.A_N(\fcounter[1] ),
    .B(FClrN),
    .X(_374_));
 sky130_fd_sc_hd__and2_2 _792_ (.A(FClrN),
    .B(\fcounter[1] ),
    .X(_375_));
 sky130_fd_sc_hd__and4bb_2 _793_ (.A_N(FOutN),
    .B_N(\fcounter[0] ),
    .C(F_EmptyN),
    .D(_348_),
    .X(_376_));
 sky130_fd_sc_hd__and4b_2 _794_ (.A_N(_348_),
    .B(_354_),
    .C(F_FullN),
    .D(FOutN),
    .X(_377_));
 sky130_fd_sc_hd__nor2_2 _795_ (.A(_376_),
    .B(_377_),
    .Y(_378_));
 sky130_fd_sc_hd__mux2_2 _796_ (.A0(_374_),
    .A1(_375_),
    .S(_378_),
    .X(_379_));
 sky130_fd_sc_hd__buf_1 _797_ (.A(_379_),
    .X(_136_));
 sky130_fd_sc_hd__and3b_2 _798_ (.A_N(_377_),
    .B(_375_),
    .C(_359_),
    .X(_380_));
 sky130_fd_sc_hd__and3b_2 _799_ (.A_N(_359_),
    .B(_377_),
    .C(_375_),
    .X(_381_));
 sky130_fd_sc_hd__and3b_2 _800_ (.A_N(_376_),
    .B(_374_),
    .C(_359_),
    .X(_382_));
 sky130_fd_sc_hd__and3b_2 _801_ (.A_N(_359_),
    .B(_376_),
    .C(_374_),
    .X(_383_));
 sky130_fd_sc_hd__or4_4 _802_ (.A(_380_),
    .B(_381_),
    .C(_382_),
    .D(_383_),
    .X(_384_));
 sky130_fd_sc_hd__buf_6 _803_ (.A(_384_),
    .X(_137_));
 sky130_fd_sc_hd__or2b_2 _804_ (.A(_352_),
    .B_N(_140_),
    .X(_385_));
 sky130_fd_sc_hd__or2_2 _805_ (.A(_347_),
    .B(_141_),
    .X(_386_));
 sky130_fd_sc_hd__and3_2 _806_ (.A(_223_),
    .B(_385_),
    .C(_386_),
    .X(_387_));
 sky130_fd_sc_hd__buf_1 _807_ (.A(_387_),
    .X(_138_));
 sky130_fd_sc_hd__xor2_2 _808_ (.A(_143_),
    .B(_385_),
    .X(_388_));
 sky130_fd_sc_hd__nor2_2 _809_ (.A(_232_),
    .B(_388_),
    .Y(_139_));
 sky130_fd_sc_hd__dfxtp_2 _810_ (.CLK(Clk),
    .D(_000_),
    .Q(\memblk.FIFO[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _811_ (.CLK(Clk),
    .D(_001_),
    .Q(\memblk.FIFO[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _812_ (.CLK(Clk),
    .D(_002_),
    .Q(\memblk.FIFO[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _813_ (.CLK(Clk),
    .D(_003_),
    .Q(\memblk.FIFO[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _814_ (.CLK(Clk),
    .D(_004_),
    .Q(\memblk.FIFO[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _815_ (.CLK(Clk),
    .D(_005_),
    .Q(\memblk.FIFO[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _816_ (.CLK(Clk),
    .D(_006_),
    .Q(\memblk.FIFO[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _817_ (.CLK(Clk),
    .D(_007_),
    .Q(\memblk.FIFO[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _818_ (.CLK(Clk),
    .D(_008_),
    .Q(\memblk.FIFO[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _819_ (.CLK(Clk),
    .D(_009_),
    .Q(\memblk.FIFO[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _820_ (.CLK(Clk),
    .D(_010_),
    .Q(\memblk.FIFO[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _821_ (.CLK(Clk),
    .D(_011_),
    .Q(\memblk.FIFO[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _822_ (.CLK(Clk),
    .D(_012_),
    .Q(\memblk.FIFO[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _823_ (.CLK(Clk),
    .D(_013_),
    .Q(\memblk.FIFO[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _824_ (.CLK(Clk),
    .D(_014_),
    .Q(\memblk.FIFO[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _825_ (.CLK(Clk),
    .D(_015_),
    .Q(\memblk.FIFO[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _826_ (.CLK(Clk),
    .D(_016_),
    .Q(\memblk.FIFO[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _827_ (.CLK(Clk),
    .D(_017_),
    .Q(\memblk.FIFO[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _828_ (.CLK(Clk),
    .D(_018_),
    .Q(\memblk.FIFO[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _829_ (.CLK(Clk),
    .D(_019_),
    .Q(\memblk.FIFO[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _830_ (.CLK(Clk),
    .D(_020_),
    .Q(\memblk.FIFO[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _831_ (.CLK(Clk),
    .D(_021_),
    .Q(\memblk.FIFO[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _832_ (.CLK(Clk),
    .D(_022_),
    .Q(\memblk.FIFO[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _833_ (.CLK(Clk),
    .D(_023_),
    .Q(\memblk.FIFO[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _834_ (.CLK(Clk),
    .D(_024_),
    .Q(\memblk.FIFO[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _835_ (.CLK(Clk),
    .D(_025_),
    .Q(\memblk.FIFO[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _836_ (.CLK(Clk),
    .D(_026_),
    .Q(\memblk.FIFO[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _837_ (.CLK(Clk),
    .D(_027_),
    .Q(\memblk.FIFO[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _838_ (.CLK(Clk),
    .D(_028_),
    .Q(\memblk.FIFO[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _839_ (.CLK(Clk),
    .D(_029_),
    .Q(\memblk.FIFO[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _840_ (.CLK(Clk),
    .D(_030_),
    .Q(\memblk.FIFO[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _841_ (.CLK(Clk),
    .D(_031_),
    .Q(\memblk.FIFO[2][31] ));
 sky130_fd_sc_hd__dfrtp_2 _842_ (.CLK(Clk),
    .D(_032_),
    .RESET_B(RstN),
    .Q(\memblk.wr_addr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _843_ (.CLK(Clk),
    .D(_033_),
    .RESET_B(RstN),
    .Q(\memblk.wr_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _844_ (.CLK(Clk),
    .D(_034_),
    .Q(\memblk.FIFO[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _845_ (.CLK(Clk),
    .D(_035_),
    .Q(\memblk.FIFO[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _846_ (.CLK(Clk),
    .D(_036_),
    .Q(\memblk.FIFO[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _847_ (.CLK(Clk),
    .D(_037_),
    .Q(\memblk.FIFO[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _848_ (.CLK(Clk),
    .D(_038_),
    .Q(\memblk.FIFO[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _849_ (.CLK(Clk),
    .D(_039_),
    .Q(\memblk.FIFO[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _850_ (.CLK(Clk),
    .D(_040_),
    .Q(\memblk.FIFO[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _851_ (.CLK(Clk),
    .D(_041_),
    .Q(\memblk.FIFO[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _852_ (.CLK(Clk),
    .D(_042_),
    .Q(\memblk.FIFO[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _853_ (.CLK(Clk),
    .D(_043_),
    .Q(\memblk.FIFO[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _854_ (.CLK(Clk),
    .D(_044_),
    .Q(\memblk.FIFO[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _855_ (.CLK(Clk),
    .D(_045_),
    .Q(\memblk.FIFO[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _856_ (.CLK(Clk),
    .D(_046_),
    .Q(\memblk.FIFO[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _857_ (.CLK(Clk),
    .D(_047_),
    .Q(\memblk.FIFO[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _858_ (.CLK(Clk),
    .D(_048_),
    .Q(\memblk.FIFO[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _859_ (.CLK(Clk),
    .D(_049_),
    .Q(\memblk.FIFO[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _860_ (.CLK(Clk),
    .D(_050_),
    .Q(\memblk.FIFO[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _861_ (.CLK(Clk),
    .D(_051_),
    .Q(\memblk.FIFO[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _862_ (.CLK(Clk),
    .D(_052_),
    .Q(\memblk.FIFO[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _863_ (.CLK(Clk),
    .D(_053_),
    .Q(\memblk.FIFO[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _864_ (.CLK(Clk),
    .D(_054_),
    .Q(\memblk.FIFO[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _865_ (.CLK(Clk),
    .D(_055_),
    .Q(\memblk.FIFO[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _866_ (.CLK(Clk),
    .D(_056_),
    .Q(\memblk.FIFO[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _867_ (.CLK(Clk),
    .D(_057_),
    .Q(\memblk.FIFO[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _868_ (.CLK(Clk),
    .D(_058_),
    .Q(\memblk.FIFO[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _869_ (.CLK(Clk),
    .D(_059_),
    .Q(\memblk.FIFO[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _870_ (.CLK(Clk),
    .D(_060_),
    .Q(\memblk.FIFO[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _871_ (.CLK(Clk),
    .D(_061_),
    .Q(\memblk.FIFO[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _872_ (.CLK(Clk),
    .D(_062_),
    .Q(\memblk.FIFO[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _873_ (.CLK(Clk),
    .D(_063_),
    .Q(\memblk.FIFO[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _874_ (.CLK(Clk),
    .D(_064_),
    .Q(\memblk.FIFO[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _875_ (.CLK(Clk),
    .D(_065_),
    .Q(\memblk.FIFO[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _876_ (.CLK(Clk),
    .D(_066_),
    .Q(\memblk.FIFO[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _877_ (.CLK(Clk),
    .D(_067_),
    .Q(\memblk.FIFO[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _878_ (.CLK(Clk),
    .D(_068_),
    .Q(\memblk.FIFO[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _879_ (.CLK(Clk),
    .D(_069_),
    .Q(\memblk.FIFO[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _880_ (.CLK(Clk),
    .D(_070_),
    .Q(\memblk.FIFO[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _881_ (.CLK(Clk),
    .D(_071_),
    .Q(\memblk.FIFO[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _882_ (.CLK(Clk),
    .D(_072_),
    .Q(\memblk.FIFO[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _883_ (.CLK(Clk),
    .D(_073_),
    .Q(\memblk.FIFO[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _884_ (.CLK(Clk),
    .D(_074_),
    .Q(\memblk.FIFO[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _885_ (.CLK(Clk),
    .D(_075_),
    .Q(\memblk.FIFO[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _886_ (.CLK(Clk),
    .D(_076_),
    .Q(\memblk.FIFO[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _887_ (.CLK(Clk),
    .D(_077_),
    .Q(\memblk.FIFO[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _888_ (.CLK(Clk),
    .D(_078_),
    .Q(\memblk.FIFO[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _889_ (.CLK(Clk),
    .D(_079_),
    .Q(\memblk.FIFO[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _890_ (.CLK(Clk),
    .D(_080_),
    .Q(\memblk.FIFO[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _891_ (.CLK(Clk),
    .D(_081_),
    .Q(\memblk.FIFO[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _892_ (.CLK(Clk),
    .D(_082_),
    .Q(\memblk.FIFO[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _893_ (.CLK(Clk),
    .D(_083_),
    .Q(\memblk.FIFO[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _894_ (.CLK(Clk),
    .D(_084_),
    .Q(\memblk.FIFO[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _895_ (.CLK(Clk),
    .D(_085_),
    .Q(\memblk.FIFO[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _896_ (.CLK(Clk),
    .D(_086_),
    .Q(\memblk.FIFO[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _897_ (.CLK(Clk),
    .D(_087_),
    .Q(\memblk.FIFO[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _898_ (.CLK(Clk),
    .D(_088_),
    .Q(\memblk.FIFO[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _899_ (.CLK(Clk),
    .D(_089_),
    .Q(\memblk.FIFO[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _900_ (.CLK(Clk),
    .D(_090_),
    .Q(\memblk.FIFO[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _901_ (.CLK(Clk),
    .D(_091_),
    .Q(\memblk.FIFO[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _902_ (.CLK(Clk),
    .D(_092_),
    .Q(\memblk.FIFO[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _903_ (.CLK(Clk),
    .D(_093_),
    .Q(\memblk.FIFO[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _904_ (.CLK(Clk),
    .D(_094_),
    .Q(\memblk.FIFO[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _905_ (.CLK(Clk),
    .D(_095_),
    .Q(\memblk.FIFO[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _906_ (.CLK(Clk),
    .D(_096_),
    .Q(\memblk.FIFO[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _907_ (.CLK(Clk),
    .D(_097_),
    .Q(\memblk.FIFO[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _908_ (.CLK(Clk),
    .D(_098_),
    .Q(\memblk.FIFO[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _909_ (.CLK(Clk),
    .D(_099_),
    .Q(\memblk.FIFO[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _910_ (.CLK(Clk),
    .D(_100_),
    .Q(\memblk.FIFO[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _911_ (.CLK(Clk),
    .D(_101_),
    .Q(\memblk.FIFO[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _912_ (.CLK(Clk),
    .D(_102_),
    .Q(\memblk.FIFO[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _913_ (.CLK(Clk),
    .D(_103_),
    .Q(\memblk.FIFO[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _914_ (.CLK(Clk),
    .D(_104_),
    .Q(\memblk.FIFO[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _915_ (.CLK(Clk),
    .D(_105_),
    .Q(\memblk.FIFO[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _916_ (.CLK(Clk),
    .D(_106_),
    .Q(\memblk.FIFO[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _917_ (.CLK(Clk),
    .D(_107_),
    .Q(\memblk.FIFO[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _918_ (.CLK(Clk),
    .D(_108_),
    .Q(\memblk.FIFO[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _919_ (.CLK(Clk),
    .D(_109_),
    .Q(\memblk.FIFO[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _920_ (.CLK(Clk),
    .D(_110_),
    .Q(\memblk.FIFO[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _921_ (.CLK(Clk),
    .D(_111_),
    .Q(\memblk.FIFO[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _922_ (.CLK(Clk),
    .D(_112_),
    .Q(\memblk.FIFO[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _923_ (.CLK(Clk),
    .D(_113_),
    .Q(\memblk.FIFO[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _924_ (.CLK(Clk),
    .D(_114_),
    .Q(\memblk.FIFO[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _925_ (.CLK(Clk),
    .D(_115_),
    .Q(\memblk.FIFO[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _926_ (.CLK(Clk),
    .D(_116_),
    .Q(\memblk.FIFO[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _927_ (.CLK(Clk),
    .D(_117_),
    .Q(\memblk.FIFO[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _928_ (.CLK(Clk),
    .D(_118_),
    .Q(\memblk.FIFO[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _929_ (.CLK(Clk),
    .D(_119_),
    .Q(\memblk.FIFO[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _930_ (.CLK(Clk),
    .D(_120_),
    .Q(\memblk.FIFO[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _931_ (.CLK(Clk),
    .D(_121_),
    .Q(\memblk.FIFO[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _932_ (.CLK(Clk),
    .D(_122_),
    .Q(\memblk.FIFO[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _933_ (.CLK(Clk),
    .D(_123_),
    .Q(\memblk.FIFO[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _934_ (.CLK(Clk),
    .D(_124_),
    .Q(\memblk.FIFO[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _935_ (.CLK(Clk),
    .D(_125_),
    .Q(\memblk.FIFO[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _936_ (.CLK(Clk),
    .D(_126_),
    .Q(\memblk.FIFO[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _937_ (.CLK(Clk),
    .D(_127_),
    .Q(\memblk.FIFO[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _938_ (.CLK(Clk),
    .D(_128_),
    .Q(\memblk.FIFO[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _939_ (.CLK(Clk),
    .D(_129_),
    .Q(\memblk.FIFO[3][31] ));
 sky130_fd_sc_hd__dfstp_2 _940_ (.CLK(Clk),
    .D(_130_),
    .SET_B(RstN),
    .Q(F_FullN));
 sky130_fd_sc_hd__dfstp_2 _941_ (.CLK(Clk),
    .D(_131_),
    .SET_B(RstN),
    .Q(F_LastN));
 sky130_fd_sc_hd__dfstp_2 _942_ (.CLK(Clk),
    .D(_132_),
    .SET_B(RstN),
    .Q(F_SLastN));
 sky130_fd_sc_hd__dfstp_2 _943_ (.CLK(Clk),
    .D(_133_),
    .SET_B(RstN),
    .Q(F_FirstN));
 sky130_fd_sc_hd__dfrtp_2 _944_ (.CLK(Clk),
    .D(_134_),
    .RESET_B(RstN),
    .Q(F_EmptyN));
 sky130_fd_sc_hd__dfrtp_2 _945_ (.CLK(Clk),
    .D(_135_),
    .RESET_B(RstN),
    .Q(\fcounter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _946_ (.CLK(Clk),
    .D(_136_),
    .RESET_B(RstN),
    .Q(\fcounter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _947_ (.CLK(Clk),
    .D(_137_),
    .RESET_B(RstN),
    .Q(\fcounter[2] ));
 sky130_fd_sc_hd__dfrtp_2 _948_ (.CLK(Clk),
    .D(_138_),
    .RESET_B(RstN),
    .Q(\memblk.rd_addr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _949_ (.CLK(Clk),
    .D(_139_),
    .RESET_B(RstN),
    .Q(\memblk.rd_addr[1] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_259 ();
endmodule
